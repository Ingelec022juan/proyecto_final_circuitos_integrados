module Timer_PWM_Generator (PWM_OUTA,
    PWM_OUTB,
    clk,
    reset,
    timer_interrupt,
    PWM_CNTA,
    PWM_CNTB,
    TIMER_TOP,
    TMR_MODE,
    TMR_SRC);
 output PWM_OUTA;
 output PWM_OUTB;
 input clk;
 input reset;
 output timer_interrupt;
 input [31:0] PWM_CNTA;
 input [31:0] PWM_CNTB;
 input [31:0] TIMER_TOP;
 input [1:0] TMR_MODE;
 input [1:0] TMR_SRC;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire \fast_pwm_inst.pwm_counter[0] ;
 wire \fast_pwm_inst.pwm_counter[10] ;
 wire \fast_pwm_inst.pwm_counter[11] ;
 wire \fast_pwm_inst.pwm_counter[12] ;
 wire \fast_pwm_inst.pwm_counter[13] ;
 wire \fast_pwm_inst.pwm_counter[14] ;
 wire \fast_pwm_inst.pwm_counter[15] ;
 wire \fast_pwm_inst.pwm_counter[16] ;
 wire \fast_pwm_inst.pwm_counter[17] ;
 wire \fast_pwm_inst.pwm_counter[18] ;
 wire \fast_pwm_inst.pwm_counter[19] ;
 wire \fast_pwm_inst.pwm_counter[1] ;
 wire \fast_pwm_inst.pwm_counter[20] ;
 wire \fast_pwm_inst.pwm_counter[21] ;
 wire \fast_pwm_inst.pwm_counter[22] ;
 wire \fast_pwm_inst.pwm_counter[23] ;
 wire \fast_pwm_inst.pwm_counter[24] ;
 wire \fast_pwm_inst.pwm_counter[25] ;
 wire \fast_pwm_inst.pwm_counter[26] ;
 wire \fast_pwm_inst.pwm_counter[27] ;
 wire \fast_pwm_inst.pwm_counter[28] ;
 wire \fast_pwm_inst.pwm_counter[29] ;
 wire \fast_pwm_inst.pwm_counter[2] ;
 wire \fast_pwm_inst.pwm_counter[30] ;
 wire \fast_pwm_inst.pwm_counter[31] ;
 wire \fast_pwm_inst.pwm_counter[3] ;
 wire \fast_pwm_inst.pwm_counter[4] ;
 wire \fast_pwm_inst.pwm_counter[5] ;
 wire \fast_pwm_inst.pwm_counter[6] ;
 wire \fast_pwm_inst.pwm_counter[7] ;
 wire \fast_pwm_inst.pwm_counter[8] ;
 wire \fast_pwm_inst.pwm_counter[9] ;
 wire \fast_pwm_inst.pwm_outa ;
 wire \fast_pwm_inst.pwm_outb ;
 wire irq_timer_normal;
 wire \normal_mode_inst.timer_cnt[0] ;
 wire \normal_mode_inst.timer_cnt[10] ;
 wire \normal_mode_inst.timer_cnt[11] ;
 wire \normal_mode_inst.timer_cnt[12] ;
 wire \normal_mode_inst.timer_cnt[13] ;
 wire \normal_mode_inst.timer_cnt[14] ;
 wire \normal_mode_inst.timer_cnt[15] ;
 wire \normal_mode_inst.timer_cnt[16] ;
 wire \normal_mode_inst.timer_cnt[17] ;
 wire \normal_mode_inst.timer_cnt[18] ;
 wire \normal_mode_inst.timer_cnt[19] ;
 wire \normal_mode_inst.timer_cnt[1] ;
 wire \normal_mode_inst.timer_cnt[20] ;
 wire \normal_mode_inst.timer_cnt[21] ;
 wire \normal_mode_inst.timer_cnt[22] ;
 wire \normal_mode_inst.timer_cnt[23] ;
 wire \normal_mode_inst.timer_cnt[24] ;
 wire \normal_mode_inst.timer_cnt[25] ;
 wire \normal_mode_inst.timer_cnt[26] ;
 wire \normal_mode_inst.timer_cnt[27] ;
 wire \normal_mode_inst.timer_cnt[28] ;
 wire \normal_mode_inst.timer_cnt[29] ;
 wire \normal_mode_inst.timer_cnt[2] ;
 wire \normal_mode_inst.timer_cnt[30] ;
 wire \normal_mode_inst.timer_cnt[31] ;
 wire \normal_mode_inst.timer_cnt[3] ;
 wire \normal_mode_inst.timer_cnt[4] ;
 wire \normal_mode_inst.timer_cnt[5] ;
 wire \normal_mode_inst.timer_cnt[6] ;
 wire \normal_mode_inst.timer_cnt[7] ;
 wire \normal_mode_inst.timer_cnt[8] ;
 wire \normal_mode_inst.timer_cnt[9] ;
 wire \phase_pwm_inst.counter[0] ;
 wire \phase_pwm_inst.counter[10] ;
 wire \phase_pwm_inst.counter[11] ;
 wire \phase_pwm_inst.counter[12] ;
 wire \phase_pwm_inst.counter[13] ;
 wire \phase_pwm_inst.counter[14] ;
 wire \phase_pwm_inst.counter[15] ;
 wire \phase_pwm_inst.counter[16] ;
 wire \phase_pwm_inst.counter[17] ;
 wire \phase_pwm_inst.counter[18] ;
 wire \phase_pwm_inst.counter[19] ;
 wire \phase_pwm_inst.counter[1] ;
 wire \phase_pwm_inst.counter[20] ;
 wire \phase_pwm_inst.counter[21] ;
 wire \phase_pwm_inst.counter[22] ;
 wire \phase_pwm_inst.counter[23] ;
 wire \phase_pwm_inst.counter[24] ;
 wire \phase_pwm_inst.counter[25] ;
 wire \phase_pwm_inst.counter[26] ;
 wire \phase_pwm_inst.counter[27] ;
 wire \phase_pwm_inst.counter[28] ;
 wire \phase_pwm_inst.counter[29] ;
 wire \phase_pwm_inst.counter[2] ;
 wire \phase_pwm_inst.counter[30] ;
 wire \phase_pwm_inst.counter[31] ;
 wire \phase_pwm_inst.counter[3] ;
 wire \phase_pwm_inst.counter[4] ;
 wire \phase_pwm_inst.counter[5] ;
 wire \phase_pwm_inst.counter[6] ;
 wire \phase_pwm_inst.counter[7] ;
 wire \phase_pwm_inst.counter[8] ;
 wire \phase_pwm_inst.counter[9] ;
 wire \phase_pwm_inst.direction ;
 wire \phase_pwm_inst.pwm_outa ;
 wire \phase_pwm_inst.pwm_outb ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__inv_2 _0942_ (.A(\phase_pwm_inst.counter[31] ),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(\phase_pwm_inst.counter[30] ),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_2 _0944_ (.A(\phase_pwm_inst.counter[29] ),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_2 _0945_ (.A(\phase_pwm_inst.counter[28] ),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_2 _0946_ (.A(\phase_pwm_inst.counter[27] ),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _0947_ (.A(\phase_pwm_inst.counter[26] ),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_2 _0948_ (.A(\phase_pwm_inst.counter[25] ),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_2 _0949_ (.A(\phase_pwm_inst.counter[24] ),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_2 _0950_ (.A(\phase_pwm_inst.counter[23] ),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_2 _0951_ (.A(\phase_pwm_inst.counter[22] ),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_2 _0952_ (.A(\phase_pwm_inst.counter[21] ),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(\phase_pwm_inst.counter[20] ),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(\phase_pwm_inst.counter[19] ),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(\phase_pwm_inst.counter[18] ),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(\phase_pwm_inst.counter[17] ),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(\phase_pwm_inst.counter[16] ),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _0958_ (.A(\phase_pwm_inst.counter[15] ),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_2 _0959_ (.A(\phase_pwm_inst.counter[14] ),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_2 _0960_ (.A(\phase_pwm_inst.counter[12] ),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _0961_ (.A(\phase_pwm_inst.counter[11] ),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(\phase_pwm_inst.counter[10] ),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _0963_ (.A(\phase_pwm_inst.counter[9] ),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_2 _0964_ (.A(\phase_pwm_inst.counter[8] ),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(\phase_pwm_inst.counter[7] ),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_2 _0966_ (.A(\phase_pwm_inst.counter[6] ),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(\phase_pwm_inst.counter[5] ),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(\phase_pwm_inst.counter[4] ),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_2 _0969_ (.A(\phase_pwm_inst.counter[3] ),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(\phase_pwm_inst.counter[2] ),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_2 _0971_ (.A(\phase_pwm_inst.counter[1] ),
    .Y(_0450_));
 sky130_fd_sc_hd__inv_2 _0972_ (.A(\phase_pwm_inst.counter[0] ),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _0973_ (.A(\normal_mode_inst.timer_cnt[0] ),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _0974_ (.A(net89),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_2 _0975_ (.A(net88),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_2 _0976_ (.A(net86),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(net85),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_2 _0978_ (.A(net84),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _0979_ (.A(net83),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(net82),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(net80),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_2 _0982_ (.A(net79),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_2 _0983_ (.A(net78),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(net72),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(net71),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_2 _0986_ (.A(net69),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_2 _0987_ (.A(net67),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_2 _0988_ (.A(net95),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_2 _0989_ (.A(net93),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(net90),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_2 _0991_ (.A(net87),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_2 _0992_ (.A(\phase_pwm_inst.direction ),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_2 _0993_ (.A(\fast_pwm_inst.pwm_counter[31] ),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(\fast_pwm_inst.pwm_counter[30] ),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_2 _0995_ (.A(\fast_pwm_inst.pwm_counter[29] ),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _0996_ (.A(\fast_pwm_inst.pwm_counter[28] ),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_2 _0997_ (.A(\fast_pwm_inst.pwm_counter[27] ),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_2 _0998_ (.A(\fast_pwm_inst.pwm_counter[26] ),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_2 _0999_ (.A(\fast_pwm_inst.pwm_counter[25] ),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(\fast_pwm_inst.pwm_counter[24] ),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(\fast_pwm_inst.pwm_counter[23] ),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_2 _1002_ (.A(\fast_pwm_inst.pwm_counter[22] ),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _1003_ (.A(\fast_pwm_inst.pwm_counter[21] ),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_2 _1004_ (.A(\fast_pwm_inst.pwm_counter[20] ),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_2 _1005_ (.A(\fast_pwm_inst.pwm_counter[19] ),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_2 _1006_ (.A(\fast_pwm_inst.pwm_counter[18] ),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _1007_ (.A(\fast_pwm_inst.pwm_counter[17] ),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _1008_ (.A(\fast_pwm_inst.pwm_counter[16] ),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_2 _1009_ (.A(\fast_pwm_inst.pwm_counter[14] ),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_2 _1010_ (.A(\fast_pwm_inst.pwm_counter[13] ),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_2 _1011_ (.A(\fast_pwm_inst.pwm_counter[12] ),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_2 _1012_ (.A(\fast_pwm_inst.pwm_counter[11] ),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _1013_ (.A(\fast_pwm_inst.pwm_counter[10] ),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_2 _1014_ (.A(\fast_pwm_inst.pwm_counter[9] ),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _1015_ (.A(\fast_pwm_inst.pwm_counter[8] ),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_2 _1016_ (.A(\fast_pwm_inst.pwm_counter[7] ),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_2 _1017_ (.A(\fast_pwm_inst.pwm_counter[6] ),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _1018_ (.A(\fast_pwm_inst.pwm_counter[5] ),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_2 _1019_ (.A(\fast_pwm_inst.pwm_counter[4] ),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_2 _1020_ (.A(\fast_pwm_inst.pwm_counter[3] ),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_2 _1021_ (.A(\fast_pwm_inst.pwm_counter[2] ),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _1022_ (.A(\fast_pwm_inst.pwm_counter[1] ),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_2 _1023_ (.A(\fast_pwm_inst.pwm_counter[0] ),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _1024_ (.A(net52),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_2 _1025_ (.A(net50),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(net49),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _1027_ (.A(net48),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(net47),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_2 _1029_ (.A(net46),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _1030_ (.A(net45),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_2 _1031_ (.A(net43),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_2 _1032_ (.A(net42),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_2 _1033_ (.A(net41),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _1034_ (.A(net40),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _1035_ (.A(net39),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(net38),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(net37),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _1038_ (.A(net36),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(net35),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _1040_ (.A(net34),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _1041_ (.A(net58),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _1042_ (.A(net22),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(net21),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _1044_ (.A(net20),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _1045_ (.A(net19),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _1046_ (.A(net18),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _1047_ (.A(net17),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _1048_ (.A(net14),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _1049_ (.A(net13),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _1050_ (.A(net11),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _1051_ (.A(net10),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _1052_ (.A(net9),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _1053_ (.A(net8),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(net7),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(net6),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(net5),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(net4),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(net2),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(net99),
    .Y(_0070_));
 sky130_fd_sc_hd__nand2_1 _1060_ (.A(_0429_),
    .B(net80),
    .Y(_0537_));
 sky130_fd_sc_hd__a22o_1 _1061_ (.A1(\phase_pwm_inst.counter[23] ),
    .A2(_0459_),
    .B1(_0460_),
    .B2(\phase_pwm_inst.counter[22] ),
    .X(_0538_));
 sky130_fd_sc_hd__o22a_1 _1062_ (.A1(\phase_pwm_inst.counter[22] ),
    .A2(_0460_),
    .B1(_0461_),
    .B2(\phase_pwm_inst.counter[21] ),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0435_),
    .B(net73),
    .Y(_0540_));
 sky130_fd_sc_hd__o22ai_1 _1064_ (.A1(_0434_),
    .A2(net74),
    .B1(net73),
    .B2(_0435_),
    .Y(_0541_));
 sky130_fd_sc_hd__a31o_1 _1065_ (.A1(\phase_pwm_inst.counter[16] ),
    .A2(_0462_),
    .A3(_0540_),
    .B1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__and2_1 _1066_ (.A(_0432_),
    .B(net77),
    .X(_0543_));
 sky130_fd_sc_hd__a21oi_1 _1067_ (.A1(_0433_),
    .A2(net75),
    .B1(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _1068_ (.A(_0434_),
    .B(net74),
    .Y(_0545_));
 sky130_fd_sc_hd__nor2_1 _1069_ (.A(_0431_),
    .B(net78),
    .Y(_0546_));
 sky130_fd_sc_hd__o22a_1 _1070_ (.A1(_0432_),
    .A2(net77),
    .B1(net75),
    .B2(_0433_),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _1071_ (.A(_0543_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a311o_1 _1072_ (.A1(_0542_),
    .A2(_0544_),
    .A3(_0545_),
    .B1(_0546_),
    .C1(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _1073_ (.A1(_0539_),
    .A2(_0549_),
    .B1(_0538_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_1 _1074_ (.A(_0438_),
    .B(net70),
    .Y(_0551_));
 sky130_fd_sc_hd__o2bb2a_1 _1075_ (.A1_N(_0439_),
    .A2_N(net68),
    .B1(_0465_),
    .B2(\phase_pwm_inst.counter[11] ),
    .X(_0552_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nand2b_1 _1077_ (.A_N(\phase_pwm_inst.counter[1] ),
    .B(net76),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2b_1 _1078_ (.A_N(\phase_pwm_inst.counter[0] ),
    .B(net65),
    .Y(_0555_));
 sky130_fd_sc_hd__and2b_1 _1079_ (.A_N(net76),
    .B(\phase_pwm_inst.counter[1] ),
    .X(_0556_));
 sky130_fd_sc_hd__a221o_1 _1080_ (.A1(\phase_pwm_inst.counter[2] ),
    .A2(_0469_),
    .B1(_0554_),
    .B2(_0555_),
    .C1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__nand2_1 _1081_ (.A(_0447_),
    .B(net91),
    .Y(_0558_));
 sky130_fd_sc_hd__o22a_1 _1082_ (.A1(\phase_pwm_inst.counter[3] ),
    .A2(_0468_),
    .B1(_0469_),
    .B2(\phase_pwm_inst.counter[2] ),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _1083_ (.A1(\phase_pwm_inst.counter[3] ),
    .A2(_0468_),
    .B1(_0557_),
    .B2(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__o22a_1 _1084_ (.A1(_0446_),
    .A2(net92),
    .B1(net91),
    .B2(_0447_),
    .X(_0561_));
 sky130_fd_sc_hd__a21bo_1 _1085_ (.A1(_0558_),
    .A2(_0560_),
    .B1_N(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__o2bb2a_1 _1086_ (.A1_N(net92),
    .A2_N(_0446_),
    .B1(\phase_pwm_inst.counter[6] ),
    .B2(_0467_),
    .X(_0563_));
 sky130_fd_sc_hd__o22a_1 _1087_ (.A1(_0444_),
    .A2(net94),
    .B1(net93),
    .B2(_0445_),
    .X(_0564_));
 sky130_fd_sc_hd__a21bo_1 _1088_ (.A1(_0562_),
    .A2(_0563_),
    .B1_N(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__o22a_1 _1089_ (.A1(_0440_),
    .A2(net67),
    .B1(net66),
    .B2(_0441_),
    .X(_0566_));
 sky130_fd_sc_hd__o221ai_2 _1090_ (.A1(_0442_),
    .A2(net96),
    .B1(net95),
    .B2(_0443_),
    .C1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__a22o_1 _1091_ (.A1(_0441_),
    .A2(net66),
    .B1(net96),
    .B2(_0442_),
    .X(_0568_));
 sky130_fd_sc_hd__nor2_1 _1092_ (.A(_0439_),
    .B(net68),
    .Y(_0569_));
 sky130_fd_sc_hd__a21oi_1 _1093_ (.A1(_0444_),
    .A2(net94),
    .B1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(\phase_pwm_inst.counter[13] ),
    .B(_0464_),
    .X(_0571_));
 sky130_fd_sc_hd__o211a_1 _1095_ (.A1(\phase_pwm_inst.counter[8] ),
    .A2(_0466_),
    .B1(_0570_),
    .C1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__a21boi_1 _1096_ (.A1(_0566_),
    .A2(_0568_),
    .B1_N(_0552_),
    .Y(_0573_));
 sky130_fd_sc_hd__a221o_1 _1097_ (.A1(\phase_pwm_inst.counter[13] ),
    .A2(_0464_),
    .B1(_0567_),
    .B2(_0573_),
    .C1(_0569_),
    .X(_0574_));
 sky130_fd_sc_hd__and2_1 _1098_ (.A(_0571_),
    .B(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nor3_1 _1099_ (.A(_0553_),
    .B(_0567_),
    .C(_0568_),
    .Y(_0576_));
 sky130_fd_sc_hd__a31o_1 _1100_ (.A1(_0565_),
    .A2(_0572_),
    .A3(_0576_),
    .B1(_0575_),
    .X(_0577_));
 sky130_fd_sc_hd__o22a_1 _1101_ (.A1(_0437_),
    .A2(net71),
    .B1(net70),
    .B2(_0438_),
    .X(_0578_));
 sky130_fd_sc_hd__a21bo_1 _1102_ (.A1(_0551_),
    .A2(_0577_),
    .B1_N(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a221oi_1 _1103_ (.A1(_0436_),
    .A2(net72),
    .B1(net71),
    .B2(_0437_),
    .C1(_0546_),
    .Y(_0580_));
 sky130_fd_sc_hd__o2111a_1 _1104_ (.A1(_0436_),
    .A2(net72),
    .B1(_0537_),
    .C1(_0540_),
    .D1(_0545_),
    .X(_0581_));
 sky130_fd_sc_hd__and4b_1 _1105_ (.A_N(_0538_),
    .B(_0539_),
    .C(_0580_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__and4b_1 _1106_ (.A_N(_0541_),
    .B(_0544_),
    .C(_0547_),
    .D(_0582_),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _1107_ (.A1(_0537_),
    .A2(_0550_),
    .B1(_0579_),
    .B2(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _1108_ (.A1(_0423_),
    .A2(net86),
    .B1(net85),
    .B2(_0424_),
    .X(_0585_));
 sky130_fd_sc_hd__nor2_1 _1109_ (.A(\phase_pwm_inst.counter[25] ),
    .B(_0458_),
    .Y(_0586_));
 sky130_fd_sc_hd__a211o_1 _1110_ (.A1(_0428_),
    .A2(net81),
    .B1(_0585_),
    .C1(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _1111_ (.A1(_0421_),
    .A2(net89),
    .B1(net88),
    .B2(_0422_),
    .X(_0588_));
 sky130_fd_sc_hd__o22a_1 _1112_ (.A1(\phase_pwm_inst.counter[27] ),
    .A2(_0456_),
    .B1(_0457_),
    .B2(\phase_pwm_inst.counter[26] ),
    .X(_0589_));
 sky130_fd_sc_hd__or3b_1 _1113_ (.A(_0587_),
    .B(_0588_),
    .C_N(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__nand2_1 _1114_ (.A(\phase_pwm_inst.counter[26] ),
    .B(_0457_),
    .Y(_0591_));
 sky130_fd_sc_hd__o221a_1 _1115_ (.A1(_0427_),
    .A2(net82),
    .B1(net81),
    .B2(_0428_),
    .C1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__o22a_1 _1116_ (.A1(_0422_),
    .A2(net88),
    .B1(net86),
    .B2(_0423_),
    .X(_0593_));
 sky130_fd_sc_hd__o221a_1 _1117_ (.A1(_0424_),
    .A2(net85),
    .B1(net84),
    .B2(_0425_),
    .C1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__and4b_1 _1118_ (.A_N(_0590_),
    .B(_0592_),
    .C(_0594_),
    .D(_0584_),
    .X(_0595_));
 sky130_fd_sc_hd__a21oi_1 _1119_ (.A1(_0586_),
    .A2(_0591_),
    .B1(_0592_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _1120_ (.A(_0589_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__a221o_1 _1121_ (.A1(_0585_),
    .A2(_0593_),
    .B1(_0594_),
    .B2(_0597_),
    .C1(_0588_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ai_1 _1122_ (.A1(_0421_),
    .A2(net89),
    .B1(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__or2_1 _1123_ (.A(_0595_),
    .B(_0599_),
    .X(_0600_));
 sky130_fd_sc_hd__or4_1 _1124_ (.A(\phase_pwm_inst.counter[3] ),
    .B(\phase_pwm_inst.counter[2] ),
    .C(\phase_pwm_inst.counter[1] ),
    .D(\phase_pwm_inst.counter[0] ),
    .X(_0601_));
 sky130_fd_sc_hd__or2_1 _1125_ (.A(\phase_pwm_inst.counter[30] ),
    .B(\phase_pwm_inst.counter[29] ),
    .X(_0602_));
 sky130_fd_sc_hd__or3_1 _1126_ (.A(\phase_pwm_inst.counter[31] ),
    .B(\phase_pwm_inst.counter[28] ),
    .C(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__or4_1 _1127_ (.A(\phase_pwm_inst.counter[7] ),
    .B(\phase_pwm_inst.counter[6] ),
    .C(\phase_pwm_inst.counter[5] ),
    .D(\phase_pwm_inst.counter[4] ),
    .X(_0604_));
 sky130_fd_sc_hd__or4_1 _1128_ (.A(\phase_pwm_inst.counter[27] ),
    .B(\phase_pwm_inst.counter[26] ),
    .C(\phase_pwm_inst.counter[25] ),
    .D(\phase_pwm_inst.counter[24] ),
    .X(_0605_));
 sky130_fd_sc_hd__or4_1 _1129_ (.A(_0601_),
    .B(_0603_),
    .C(_0604_),
    .D(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__or4_1 _1130_ (.A(\phase_pwm_inst.counter[19] ),
    .B(\phase_pwm_inst.counter[18] ),
    .C(\phase_pwm_inst.counter[17] ),
    .D(\phase_pwm_inst.counter[16] ),
    .X(_0607_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(\phase_pwm_inst.direction ),
    .B(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__or4_1 _1132_ (.A(\phase_pwm_inst.counter[23] ),
    .B(\phase_pwm_inst.counter[22] ),
    .C(\phase_pwm_inst.counter[21] ),
    .D(\phase_pwm_inst.counter[20] ),
    .X(_0609_));
 sky130_fd_sc_hd__or2_1 _1133_ (.A(_0607_),
    .B(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__or4_1 _1134_ (.A(\phase_pwm_inst.counter[11] ),
    .B(\phase_pwm_inst.counter[10] ),
    .C(\phase_pwm_inst.counter[9] ),
    .D(\phase_pwm_inst.counter[8] ),
    .X(_0611_));
 sky130_fd_sc_hd__and2_1 _1135_ (.A(\phase_pwm_inst.direction ),
    .B(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__or4_1 _1136_ (.A(\phase_pwm_inst.counter[15] ),
    .B(\phase_pwm_inst.counter[14] ),
    .C(\phase_pwm_inst.counter[13] ),
    .D(\phase_pwm_inst.counter[12] ),
    .X(_0613_));
 sky130_fd_sc_hd__or2_1 _1137_ (.A(_0611_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__o31a_1 _1138_ (.A1(_0606_),
    .A2(_0610_),
    .A3(_0614_),
    .B1(\phase_pwm_inst.direction ),
    .X(_0615_));
 sky130_fd_sc_hd__o21ba_4 _1139_ (.A1(\phase_pwm_inst.direction ),
    .A2(_0600_),
    .B1_N(_0615_),
    .X(_0616_));
 sky130_fd_sc_hd__nor2_1 _1140_ (.A(_0447_),
    .B(_0470_),
    .Y(_0617_));
 sky130_fd_sc_hd__nor2_1 _1141_ (.A(\phase_pwm_inst.counter[4] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0618_));
 sky130_fd_sc_hd__nor2_1 _1142_ (.A(_0617_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__nor2_1 _1143_ (.A(\phase_pwm_inst.counter[3] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0620_));
 sky130_fd_sc_hd__or2_1 _1144_ (.A(\phase_pwm_inst.counter[3] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0621_));
 sky130_fd_sc_hd__nor2_1 _1145_ (.A(_0448_),
    .B(_0470_),
    .Y(_0622_));
 sky130_fd_sc_hd__and2_1 _1146_ (.A(\phase_pwm_inst.counter[2] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0623_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(\phase_pwm_inst.counter[1] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0624_));
 sky130_fd_sc_hd__or2_1 _1148_ (.A(\phase_pwm_inst.counter[1] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0625_));
 sky130_fd_sc_hd__nand2_1 _1149_ (.A(_0624_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__a21bo_1 _1150_ (.A1(\phase_pwm_inst.counter[0] ),
    .A2(_0625_),
    .B1_N(_0624_),
    .X(_0627_));
 sky130_fd_sc_hd__nor2_1 _1151_ (.A(\phase_pwm_inst.counter[2] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0628_));
 sky130_fd_sc_hd__nor2_1 _1152_ (.A(_0623_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a21oi_1 _1153_ (.A1(_0627_),
    .A2(_0629_),
    .B1(_0623_),
    .Y(_0630_));
 sky130_fd_sc_hd__a211o_1 _1154_ (.A1(_0627_),
    .A2(_0629_),
    .B1(_0622_),
    .C1(_0623_),
    .X(_0631_));
 sky130_fd_sc_hd__and3_1 _1155_ (.A(_0619_),
    .B(_0621_),
    .C(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_1 _1156_ (.A(_0446_),
    .B(_0470_),
    .Y(_0633_));
 sky130_fd_sc_hd__nor2_1 _1157_ (.A(\phase_pwm_inst.counter[5] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0634_));
 sky130_fd_sc_hd__nor2_1 _1158_ (.A(_0633_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__xor2_1 _1159_ (.A(\phase_pwm_inst.counter[7] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0636_));
 sky130_fd_sc_hd__nor2_1 _1160_ (.A(_0445_),
    .B(_0470_),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_1 _1161_ (.A(\phase_pwm_inst.counter[6] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0638_));
 sky130_fd_sc_hd__nor2_1 _1162_ (.A(_0637_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__and3_1 _1163_ (.A(_0635_),
    .B(_0636_),
    .C(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _1164_ (.A1(\phase_pwm_inst.direction ),
    .A2(_0604_),
    .B1(_0632_),
    .B2(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__xor2_1 _1165_ (.A(\phase_pwm_inst.counter[8] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0642_));
 sky130_fd_sc_hd__and2_1 _1166_ (.A(_0641_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__xor2_1 _1167_ (.A(\phase_pwm_inst.counter[10] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_1 _1168_ (.A(_0442_),
    .B(_0470_),
    .Y(_0645_));
 sky130_fd_sc_hd__or2_1 _1169_ (.A(\phase_pwm_inst.counter[9] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0646_));
 sky130_fd_sc_hd__nand2b_1 _1170_ (.A_N(_0645_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__xor2_1 _1171_ (.A(\phase_pwm_inst.counter[11] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0648_));
 sky130_fd_sc_hd__and4b_1 _1172_ (.A_N(_0645_),
    .B(_0646_),
    .C(_0648_),
    .D(_0644_),
    .X(_0649_));
 sky130_fd_sc_hd__and3_1 _1173_ (.A(_0641_),
    .B(_0642_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__and2_1 _1174_ (.A(\phase_pwm_inst.counter[13] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0651_));
 sky130_fd_sc_hd__or2_1 _1175_ (.A(\phase_pwm_inst.counter[13] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0652_));
 sky130_fd_sc_hd__and2b_1 _1176_ (.A_N(_0651_),
    .B(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__xor2_1 _1177_ (.A(\phase_pwm_inst.counter[14] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0654_));
 sky130_fd_sc_hd__xor2_1 _1178_ (.A(\phase_pwm_inst.counter[12] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0655_));
 sky130_fd_sc_hd__xnor2_1 _1179_ (.A(\phase_pwm_inst.counter[15] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0656_));
 sky130_fd_sc_hd__and4b_1 _1180_ (.A_N(_0656_),
    .B(_0655_),
    .C(_0654_),
    .D(_0653_),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _1181_ (.A1(\phase_pwm_inst.direction ),
    .A2(_0614_),
    .B1(_0650_),
    .B2(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__or2_1 _1182_ (.A(\phase_pwm_inst.counter[16] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0659_));
 sky130_fd_sc_hd__nand2_1 _1183_ (.A(\phase_pwm_inst.counter[16] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _1184_ (.A(_0659_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nand2b_1 _1185_ (.A_N(_0661_),
    .B(_0658_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand2_1 _1186_ (.A(\phase_pwm_inst.counter[17] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0663_));
 sky130_fd_sc_hd__nor2_1 _1187_ (.A(\phase_pwm_inst.counter[17] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _1188_ (.A(\phase_pwm_inst.counter[17] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(_0663_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__xor2_1 _1190_ (.A(\phase_pwm_inst.counter[19] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0667_));
 sky130_fd_sc_hd__xnor2_1 _1191_ (.A(\phase_pwm_inst.counter[18] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0668_));
 sky130_fd_sc_hd__and4b_1 _1192_ (.A_N(_0668_),
    .B(_0667_),
    .C(_0665_),
    .D(_0663_),
    .X(_0669_));
 sky130_fd_sc_hd__nand3b_1 _1193_ (.A_N(_0661_),
    .B(_0669_),
    .C(_0658_),
    .Y(_0670_));
 sky130_fd_sc_hd__xor2_1 _1194_ (.A(\phase_pwm_inst.counter[20] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0671_));
 sky130_fd_sc_hd__xor2_1 _1195_ (.A(\phase_pwm_inst.counter[23] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0672_));
 sky130_fd_sc_hd__nand2_1 _1196_ (.A(_0671_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__nor2_1 _1197_ (.A(_0431_),
    .B(_0470_),
    .Y(_0674_));
 sky130_fd_sc_hd__or2_1 _1198_ (.A(\phase_pwm_inst.counter[21] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0675_));
 sky130_fd_sc_hd__nand2b_1 _1199_ (.A_N(_0674_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__xnor2_2 _1200_ (.A(\phase_pwm_inst.counter[22] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0677_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__or3_1 _1202_ (.A(_0673_),
    .B(_0676_),
    .C(_0677_),
    .X(_0679_));
 sky130_fd_sc_hd__o2bb2a_1 _1203_ (.A1_N(\phase_pwm_inst.direction ),
    .A2_N(_0610_),
    .B1(_0670_),
    .B2(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__or2_1 _1204_ (.A(\phase_pwm_inst.counter[26] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(\phase_pwm_inst.counter[26] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(_0681_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__xnor2_1 _1207_ (.A(\phase_pwm_inst.counter[27] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _1208_ (.A(\phase_pwm_inst.counter[25] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0685_));
 sky130_fd_sc_hd__inv_2 _1209_ (.A(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_1 _1210_ (.A(\phase_pwm_inst.counter[25] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_1 _1211_ (.A(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nor2_1 _1212_ (.A(\phase_pwm_inst.counter[24] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1213_ (.A(\phase_pwm_inst.counter[24] ),
    .B(\phase_pwm_inst.direction ),
    .Y(_0690_));
 sky130_fd_sc_hd__and2b_1 _1214_ (.A_N(_0689_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__or4bb_1 _1215_ (.A(_0683_),
    .B(_0684_),
    .C_N(_0688_),
    .D_N(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__o2bb2a_1 _1216_ (.A1_N(\phase_pwm_inst.direction ),
    .A2_N(_0605_),
    .B1(_0680_),
    .B2(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__xor2_1 _1217_ (.A(\phase_pwm_inst.counter[28] ),
    .B(\phase_pwm_inst.direction ),
    .X(_0694_));
 sky130_fd_sc_hd__or3b_1 _1218_ (.A(\phase_pwm_inst.counter[28] ),
    .B(_0470_),
    .C_N(_0693_),
    .X(_0695_));
 sky130_fd_sc_hd__or4_1 _1219_ (.A(_0424_),
    .B(\phase_pwm_inst.direction ),
    .C(_0680_),
    .D(_0692_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _1220_ (.A(\phase_pwm_inst.counter[30] ),
    .B(\phase_pwm_inst.counter[29] ),
    .Y(_0697_));
 sky130_fd_sc_hd__a221o_1 _1221_ (.A1(_0602_),
    .A2(_0696_),
    .B1(_0697_),
    .B2(_0695_),
    .C1(_0616_),
    .X(_0698_));
 sky130_fd_sc_hd__xnor2_1 _1222_ (.A(\phase_pwm_inst.counter[31] ),
    .B(_0698_),
    .Y(_0203_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(\phase_pwm_inst.counter[29] ),
    .B(_0696_),
    .X(_0699_));
 sky130_fd_sc_hd__a211o_1 _1224_ (.A1(_0423_),
    .A2(_0695_),
    .B1(_0699_),
    .C1(_0616_),
    .X(_0700_));
 sky130_fd_sc_hd__xnor2_1 _1225_ (.A(\phase_pwm_inst.counter[30] ),
    .B(_0700_),
    .Y(_0202_));
 sky130_fd_sc_hd__a21oi_1 _1226_ (.A1(_0695_),
    .A2(_0696_),
    .B1(_0616_),
    .Y(_0701_));
 sky130_fd_sc_hd__xnor2_1 _1227_ (.A(_0423_),
    .B(_0701_),
    .Y(_0201_));
 sky130_fd_sc_hd__xnor2_1 _1228_ (.A(_0693_),
    .B(_0694_),
    .Y(_0702_));
 sky130_fd_sc_hd__mux2_1 _1229_ (.A0(_0702_),
    .A1(\phase_pwm_inst.counter[28] ),
    .S(_0616_),
    .X(_0200_));
 sky130_fd_sc_hd__o21a_1 _1230_ (.A1(_0680_),
    .A2(_0689_),
    .B1(_0690_),
    .X(_0703_));
 sky130_fd_sc_hd__o211a_1 _1231_ (.A1(_0680_),
    .A2(_0689_),
    .B1(_0690_),
    .C1(_0685_),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _1232_ (.A(_0687_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__o31a_1 _1233_ (.A1(_0683_),
    .A2(_0687_),
    .A3(_0704_),
    .B1(_0682_),
    .X(_0706_));
 sky130_fd_sc_hd__xor2_1 _1234_ (.A(_0684_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _1235_ (.A0(_0707_),
    .A1(\phase_pwm_inst.counter[27] ),
    .S(_0616_),
    .X(_0199_));
 sky130_fd_sc_hd__xnor2_1 _1236_ (.A(_0683_),
    .B(_0705_),
    .Y(_0708_));
 sky130_fd_sc_hd__mux2_1 _1237_ (.A0(_0708_),
    .A1(\phase_pwm_inst.counter[26] ),
    .S(_0616_),
    .X(_0198_));
 sky130_fd_sc_hd__xnor2_1 _1238_ (.A(_0688_),
    .B(_0703_),
    .Y(_0709_));
 sky130_fd_sc_hd__mux2_1 _1239_ (.A0(_0709_),
    .A1(\phase_pwm_inst.counter[25] ),
    .S(_0616_),
    .X(_0197_));
 sky130_fd_sc_hd__xnor2_1 _1240_ (.A(_0680_),
    .B(_0691_),
    .Y(_0710_));
 sky130_fd_sc_hd__mux2_1 _1241_ (.A0(_0710_),
    .A1(\phase_pwm_inst.counter[24] ),
    .S(_0616_),
    .X(_0196_));
 sky130_fd_sc_hd__nand2_1 _1242_ (.A(_0608_),
    .B(_0670_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21boi_1 _1243_ (.A1(_0608_),
    .A2(_0670_),
    .B1_N(_0671_),
    .Y(_0712_));
 sky130_fd_sc_hd__a21o_1 _1244_ (.A1(\phase_pwm_inst.counter[20] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a211o_1 _1245_ (.A1(\phase_pwm_inst.counter[20] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0674_),
    .C1(_0712_),
    .X(_0714_));
 sky130_fd_sc_hd__nand2_1 _1246_ (.A(_0675_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__a32o_1 _1247_ (.A1(_0675_),
    .A2(_0678_),
    .A3(_0714_),
    .B1(\phase_pwm_inst.direction ),
    .B2(\phase_pwm_inst.counter[22] ),
    .X(_0716_));
 sky130_fd_sc_hd__xor2_1 _1248_ (.A(_0672_),
    .B(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(_0717_),
    .A1(\phase_pwm_inst.counter[23] ),
    .S(_0616_),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(_0677_),
    .B(_0715_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21ba_1 _1251_ (.A1(_0677_),
    .A2(_0715_),
    .B1_N(_0616_),
    .X(_0719_));
 sky130_fd_sc_hd__a22o_1 _1252_ (.A1(\phase_pwm_inst.counter[22] ),
    .A2(_0616_),
    .B1(_0718_),
    .B2(_0719_),
    .X(_0194_));
 sky130_fd_sc_hd__xnor2_1 _1253_ (.A(_0676_),
    .B(_0713_),
    .Y(_0720_));
 sky130_fd_sc_hd__mux2_1 _1254_ (.A0(_0720_),
    .A1(\phase_pwm_inst.counter[21] ),
    .S(_0616_),
    .X(_0193_));
 sky130_fd_sc_hd__xor2_1 _1255_ (.A(_0671_),
    .B(_0711_),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1256_ (.A0(_0721_),
    .A1(\phase_pwm_inst.counter[20] ),
    .S(_0616_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(_0660_),
    .B(_0662_),
    .Y(_0722_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0665_),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a311oi_1 _1259_ (.A1(_0660_),
    .A2(_0662_),
    .A3(_0663_),
    .B1(_0664_),
    .C1(_0668_),
    .Y(_0724_));
 sky130_fd_sc_hd__a21oi_1 _1260_ (.A1(\phase_pwm_inst.counter[18] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__xnor2_1 _1261_ (.A(_0667_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__mux2_1 _1262_ (.A0(_0726_),
    .A1(\phase_pwm_inst.counter[19] ),
    .S(_0616_),
    .X(_0191_));
 sky130_fd_sc_hd__a31o_1 _1263_ (.A1(_0663_),
    .A2(_0668_),
    .A3(_0723_),
    .B1(_0616_),
    .X(_0727_));
 sky130_fd_sc_hd__a2bb2o_1 _1264_ (.A1_N(_0724_),
    .A2_N(_0727_),
    .B1(\phase_pwm_inst.counter[18] ),
    .B2(_0616_),
    .X(_0190_));
 sky130_fd_sc_hd__xnor2_1 _1265_ (.A(_0666_),
    .B(_0722_),
    .Y(_0728_));
 sky130_fd_sc_hd__mux2_1 _1266_ (.A0(_0728_),
    .A1(\phase_pwm_inst.counter[17] ),
    .S(_0616_),
    .X(_0189_));
 sky130_fd_sc_hd__and2b_1 _1267_ (.A_N(_0658_),
    .B(_0661_),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _1268_ (.A(_0616_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__a22o_1 _1269_ (.A1(\phase_pwm_inst.counter[16] ),
    .A2(_0616_),
    .B1(_0662_),
    .B2(_0730_),
    .X(_0188_));
 sky130_fd_sc_hd__o21a_1 _1270_ (.A1(_0612_),
    .A2(_0650_),
    .B1(_0655_),
    .X(_0731_));
 sky130_fd_sc_hd__a21o_1 _1271_ (.A1(\phase_pwm_inst.counter[12] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__or2_1 _1272_ (.A(_0651_),
    .B(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__nand2_1 _1273_ (.A(_0652_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__a32o_1 _1274_ (.A1(_0652_),
    .A2(_0654_),
    .A3(_0733_),
    .B1(\phase_pwm_inst.direction ),
    .B2(\phase_pwm_inst.counter[14] ),
    .X(_0735_));
 sky130_fd_sc_hd__xnor2_1 _1275_ (.A(_0656_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(_0736_),
    .A1(\phase_pwm_inst.counter[15] ),
    .S(_0616_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _1277_ (.A(_0654_),
    .B(_0734_),
    .Y(_0737_));
 sky130_fd_sc_hd__mux2_1 _1278_ (.A0(_0737_),
    .A1(\phase_pwm_inst.counter[14] ),
    .S(_0616_),
    .X(_0186_));
 sky130_fd_sc_hd__xor2_1 _1279_ (.A(_0653_),
    .B(_0732_),
    .X(_0738_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(_0738_),
    .A1(\phase_pwm_inst.counter[13] ),
    .S(_0616_),
    .X(_0185_));
 sky130_fd_sc_hd__nor3_1 _1281_ (.A(_0612_),
    .B(_0650_),
    .C(_0655_),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_1 _1282_ (.A(_0731_),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__mux2_1 _1283_ (.A0(_0740_),
    .A1(\phase_pwm_inst.counter[12] ),
    .S(_0616_),
    .X(_0184_));
 sky130_fd_sc_hd__a21o_1 _1284_ (.A1(\phase_pwm_inst.counter[8] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0643_),
    .X(_0741_));
 sky130_fd_sc_hd__o21ai_1 _1285_ (.A1(_0645_),
    .A2(_0741_),
    .B1(_0646_),
    .Y(_0742_));
 sky130_fd_sc_hd__and2b_1 _1286_ (.A_N(_0742_),
    .B(_0644_),
    .X(_0743_));
 sky130_fd_sc_hd__a21oi_1 _1287_ (.A1(\phase_pwm_inst.counter[10] ),
    .A2(\phase_pwm_inst.direction ),
    .B1(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_1 _1288_ (.A(_0648_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__mux2_1 _1289_ (.A0(_0745_),
    .A1(\phase_pwm_inst.counter[11] ),
    .S(_0616_),
    .X(_0183_));
 sky130_fd_sc_hd__xnor2_1 _1290_ (.A(_0644_),
    .B(_0742_),
    .Y(_0746_));
 sky130_fd_sc_hd__mux2_1 _1291_ (.A0(_0746_),
    .A1(\phase_pwm_inst.counter[10] ),
    .S(_0616_),
    .X(_0182_));
 sky130_fd_sc_hd__xnor2_1 _1292_ (.A(_0647_),
    .B(_0741_),
    .Y(_0747_));
 sky130_fd_sc_hd__mux2_1 _1293_ (.A0(_0747_),
    .A1(\phase_pwm_inst.counter[9] ),
    .S(_0616_),
    .X(_0181_));
 sky130_fd_sc_hd__o21bai_1 _1294_ (.A1(_0641_),
    .A2(_0642_),
    .B1_N(_0616_),
    .Y(_0748_));
 sky130_fd_sc_hd__a2bb2o_1 _1295_ (.A1_N(_0643_),
    .A2_N(_0748_),
    .B1(\phase_pwm_inst.counter[8] ),
    .B2(_0616_),
    .X(_0180_));
 sky130_fd_sc_hd__nor2_1 _1296_ (.A(_0617_),
    .B(_0632_),
    .Y(_0749_));
 sky130_fd_sc_hd__nor2_1 _1297_ (.A(_0634_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _1298_ (.A(_0633_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__o21ba_1 _1299_ (.A1(_0638_),
    .A2(_0751_),
    .B1_N(_0637_),
    .X(_0752_));
 sky130_fd_sc_hd__xnor2_1 _1300_ (.A(_0636_),
    .B(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__mux2_1 _1301_ (.A0(_0753_),
    .A1(\phase_pwm_inst.counter[7] ),
    .S(_0616_),
    .X(_0179_));
 sky130_fd_sc_hd__xnor2_1 _1302_ (.A(_0639_),
    .B(_0751_),
    .Y(_0754_));
 sky130_fd_sc_hd__mux2_1 _1303_ (.A0(_0754_),
    .A1(\phase_pwm_inst.counter[6] ),
    .S(_0616_),
    .X(_0178_));
 sky130_fd_sc_hd__xnor2_1 _1304_ (.A(_0635_),
    .B(_0749_),
    .Y(_0755_));
 sky130_fd_sc_hd__mux2_1 _1305_ (.A0(_0755_),
    .A1(\phase_pwm_inst.counter[5] ),
    .S(_0616_),
    .X(_0177_));
 sky130_fd_sc_hd__a21o_1 _1306_ (.A1(_0621_),
    .A2(_0631_),
    .B1(_0619_),
    .X(_0756_));
 sky130_fd_sc_hd__and2b_1 _1307_ (.A_N(_0632_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _1308_ (.A0(_0757_),
    .A1(\phase_pwm_inst.counter[4] ),
    .S(_0616_),
    .X(_0176_));
 sky130_fd_sc_hd__nor2_1 _1309_ (.A(_0620_),
    .B(_0622_),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _1310_ (.A(_0630_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__mux2_1 _1311_ (.A0(_0759_),
    .A1(\phase_pwm_inst.counter[3] ),
    .S(_0616_),
    .X(_0175_));
 sky130_fd_sc_hd__xor2_1 _1312_ (.A(_0627_),
    .B(_0629_),
    .X(_0760_));
 sky130_fd_sc_hd__mux2_1 _1313_ (.A0(_0760_),
    .A1(\phase_pwm_inst.counter[2] ),
    .S(_0616_),
    .X(_0174_));
 sky130_fd_sc_hd__xnor2_1 _1314_ (.A(\phase_pwm_inst.counter[0] ),
    .B(_0626_),
    .Y(_0761_));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(_0761_),
    .A1(\phase_pwm_inst.counter[1] ),
    .S(_0616_),
    .X(_0173_));
 sky130_fd_sc_hd__xnor2_1 _1316_ (.A(\phase_pwm_inst.counter[0] ),
    .B(_0616_),
    .Y(_0172_));
 sky130_fd_sc_hd__and3_1 _1317_ (.A(\normal_mode_inst.timer_cnt[0] ),
    .B(\normal_mode_inst.timer_cnt[1] ),
    .C(\normal_mode_inst.timer_cnt[2] ),
    .X(_0762_));
 sky130_fd_sc_hd__and4_1 _1318_ (.A(\normal_mode_inst.timer_cnt[0] ),
    .B(\normal_mode_inst.timer_cnt[1] ),
    .C(\normal_mode_inst.timer_cnt[3] ),
    .D(\normal_mode_inst.timer_cnt[2] ),
    .X(_0763_));
 sky130_fd_sc_hd__nand2_1 _1319_ (.A(\normal_mode_inst.timer_cnt[4] ),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__and4_1 _1320_ (.A(\normal_mode_inst.timer_cnt[5] ),
    .B(\normal_mode_inst.timer_cnt[4] ),
    .C(\normal_mode_inst.timer_cnt[6] ),
    .D(_0763_),
    .X(_0765_));
 sky130_fd_sc_hd__nand2_1 _1321_ (.A(\normal_mode_inst.timer_cnt[7] ),
    .B(_0765_),
    .Y(_0766_));
 sky130_fd_sc_hd__and4_1 _1322_ (.A(\normal_mode_inst.timer_cnt[7] ),
    .B(\normal_mode_inst.timer_cnt[9] ),
    .C(\normal_mode_inst.timer_cnt[8] ),
    .D(_0765_),
    .X(_0767_));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(\normal_mode_inst.timer_cnt[10] ),
    .B(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__and4_1 _1324_ (.A(\normal_mode_inst.timer_cnt[11] ),
    .B(\normal_mode_inst.timer_cnt[10] ),
    .C(\normal_mode_inst.timer_cnt[12] ),
    .D(_0767_),
    .X(_0769_));
 sky130_fd_sc_hd__nand2_1 _1325_ (.A(\normal_mode_inst.timer_cnt[13] ),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__and4_1 _1326_ (.A(\normal_mode_inst.timer_cnt[13] ),
    .B(\normal_mode_inst.timer_cnt[15] ),
    .C(\normal_mode_inst.timer_cnt[14] ),
    .D(_0769_),
    .X(_0771_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(\normal_mode_inst.timer_cnt[16] ),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__and4_1 _1328_ (.A(\normal_mode_inst.timer_cnt[17] ),
    .B(\normal_mode_inst.timer_cnt[16] ),
    .C(\normal_mode_inst.timer_cnt[18] ),
    .D(_0771_),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_1 _1329_ (.A(\normal_mode_inst.timer_cnt[19] ),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__and4_1 _1330_ (.A(\normal_mode_inst.timer_cnt[19] ),
    .B(\normal_mode_inst.timer_cnt[21] ),
    .C(\normal_mode_inst.timer_cnt[20] ),
    .D(_0773_),
    .X(_0775_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(\normal_mode_inst.timer_cnt[22] ),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__and4_1 _1332_ (.A(\normal_mode_inst.timer_cnt[23] ),
    .B(\normal_mode_inst.timer_cnt[22] ),
    .C(\normal_mode_inst.timer_cnt[24] ),
    .D(_0775_),
    .X(_0777_));
 sky130_fd_sc_hd__and3_1 _1333_ (.A(\normal_mode_inst.timer_cnt[25] ),
    .B(\normal_mode_inst.timer_cnt[26] ),
    .C(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__and2_1 _1334_ (.A(\normal_mode_inst.timer_cnt[27] ),
    .B(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__and3_1 _1335_ (.A(\normal_mode_inst.timer_cnt[29] ),
    .B(\normal_mode_inst.timer_cnt[28] ),
    .C(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__and3_1 _1336_ (.A(\normal_mode_inst.timer_cnt[30] ),
    .B(\normal_mode_inst.timer_cnt[31] ),
    .C(_0780_),
    .X(_0034_));
 sky130_fd_sc_hd__o22a_1 _1337_ (.A1(_0453_),
    .A2(\fast_pwm_inst.pwm_counter[30] ),
    .B1(\fast_pwm_inst.pwm_counter[29] ),
    .B2(_0454_),
    .X(_0781_));
 sky130_fd_sc_hd__o22a_1 _1338_ (.A1(_0456_),
    .A2(\fast_pwm_inst.pwm_counter[27] ),
    .B1(\fast_pwm_inst.pwm_counter[26] ),
    .B2(_0457_),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _1339_ (.A1(_0457_),
    .A2(\fast_pwm_inst.pwm_counter[26] ),
    .B1(\fast_pwm_inst.pwm_counter[25] ),
    .B2(_0458_),
    .X(_0783_));
 sky130_fd_sc_hd__a211oi_1 _1340_ (.A1(net82),
    .A2(_0477_),
    .B1(_0478_),
    .C1(net81),
    .Y(_0784_));
 sky130_fd_sc_hd__o21a_1 _1341_ (.A1(_0783_),
    .A2(_0784_),
    .B1(_0782_),
    .X(_0785_));
 sky130_fd_sc_hd__nor2_1 _1342_ (.A(net84),
    .B(_0475_),
    .Y(_0786_));
 sky130_fd_sc_hd__o22a_1 _1343_ (.A1(_0455_),
    .A2(\fast_pwm_inst.pwm_counter[28] ),
    .B1(_0785_),
    .B2(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__a221o_1 _1344_ (.A1(_0454_),
    .A2(\fast_pwm_inst.pwm_counter[29] ),
    .B1(\fast_pwm_inst.pwm_counter[28] ),
    .B2(_0455_),
    .C1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _1345_ (.A1(_0452_),
    .A2(\fast_pwm_inst.pwm_counter[31] ),
    .B1(\fast_pwm_inst.pwm_counter[30] ),
    .B2(_0453_),
    .X(_0789_));
 sky130_fd_sc_hd__a21oi_1 _1346_ (.A1(_0781_),
    .A2(_0788_),
    .B1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nor2_1 _1347_ (.A(_0452_),
    .B(\fast_pwm_inst.pwm_counter[31] ),
    .Y(_0791_));
 sky130_fd_sc_hd__nor2_1 _1348_ (.A(_0459_),
    .B(\fast_pwm_inst.pwm_counter[23] ),
    .Y(_0792_));
 sky130_fd_sc_hd__a22o_1 _1349_ (.A1(_0459_),
    .A2(\fast_pwm_inst.pwm_counter[23] ),
    .B1(\fast_pwm_inst.pwm_counter[22] ),
    .B2(_0460_),
    .X(_0793_));
 sky130_fd_sc_hd__o22a_1 _1350_ (.A1(_0460_),
    .A2(\fast_pwm_inst.pwm_counter[22] ),
    .B1(\fast_pwm_inst.pwm_counter[21] ),
    .B2(_0461_),
    .X(_0794_));
 sky130_fd_sc_hd__and2_1 _1351_ (.A(net77),
    .B(_0482_),
    .X(_0795_));
 sky130_fd_sc_hd__o22a_1 _1352_ (.A1(net73),
    .A2(_0485_),
    .B1(_0486_),
    .B2(net72),
    .X(_0796_));
 sky130_fd_sc_hd__o22a_1 _1353_ (.A1(net75),
    .A2(_0483_),
    .B1(_0484_),
    .B2(net74),
    .X(_0797_));
 sky130_fd_sc_hd__and2_1 _1354_ (.A(net75),
    .B(_0483_),
    .X(_0798_));
 sky130_fd_sc_hd__a22o_1 _1355_ (.A1(net74),
    .A2(_0484_),
    .B1(_0485_),
    .B2(net73),
    .X(_0799_));
 sky130_fd_sc_hd__or3b_1 _1356_ (.A(_0798_),
    .B(_0799_),
    .C_N(_0797_),
    .X(_0800_));
 sky130_fd_sc_hd__or2_1 _1357_ (.A(net77),
    .B(_0482_),
    .X(_0801_));
 sky130_fd_sc_hd__o221a_1 _1358_ (.A1(_0797_),
    .A2(_0798_),
    .B1(_0800_),
    .B2(_0796_),
    .C1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__a2bb2o_1 _1359_ (.A1_N(_0795_),
    .A2_N(_0802_),
    .B1(_0461_),
    .B2(\fast_pwm_inst.pwm_counter[21] ),
    .X(_0803_));
 sky130_fd_sc_hd__a21oi_1 _1360_ (.A1(_0794_),
    .A2(_0803_),
    .B1(_0793_),
    .Y(_0804_));
 sky130_fd_sc_hd__and2_1 _1361_ (.A(net91),
    .B(_0497_),
    .X(_0805_));
 sky130_fd_sc_hd__nand2b_1 _1362_ (.A_N(\fast_pwm_inst.pwm_counter[1] ),
    .B(net76),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2b_1 _1363_ (.A_N(\fast_pwm_inst.pwm_counter[0] ),
    .B(net65),
    .Y(_0807_));
 sky130_fd_sc_hd__and2b_1 _1364_ (.A_N(net76),
    .B(\fast_pwm_inst.pwm_counter[1] ),
    .X(_0808_));
 sky130_fd_sc_hd__a221o_1 _1365_ (.A1(_0469_),
    .A2(\fast_pwm_inst.pwm_counter[2] ),
    .B1(_0806_),
    .B2(_0807_),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__o22a_1 _1366_ (.A1(_0468_),
    .A2(\fast_pwm_inst.pwm_counter[3] ),
    .B1(\fast_pwm_inst.pwm_counter[2] ),
    .B2(_0469_),
    .X(_0810_));
 sky130_fd_sc_hd__o22a_1 _1367_ (.A1(net91),
    .A2(_0497_),
    .B1(_0498_),
    .B2(net90),
    .X(_0811_));
 sky130_fd_sc_hd__a21boi_1 _1368_ (.A1(_0809_),
    .A2(_0810_),
    .B1_N(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__o22a_1 _1369_ (.A1(net92),
    .A2(_0496_),
    .B1(_0805_),
    .B2(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__a22o_1 _1370_ (.A1(net93),
    .A2(_0495_),
    .B1(_0496_),
    .B2(net92),
    .X(_0814_));
 sky130_fd_sc_hd__nand2_1 _1371_ (.A(_0467_),
    .B(\fast_pwm_inst.pwm_counter[6] ),
    .Y(_0815_));
 sky130_fd_sc_hd__o221a_1 _1372_ (.A1(net94),
    .A2(_0494_),
    .B1(_0813_),
    .B2(_0814_),
    .C1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__and2_1 _1373_ (.A(net96),
    .B(_0492_),
    .X(_0817_));
 sky130_fd_sc_hd__a221o_1 _1374_ (.A1(net95),
    .A2(_0493_),
    .B1(_0494_),
    .B2(net94),
    .C1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__nand2_1 _1375_ (.A(_0466_),
    .B(\fast_pwm_inst.pwm_counter[8] ),
    .Y(_0819_));
 sky130_fd_sc_hd__o221a_1 _1376_ (.A1(net96),
    .A2(_0492_),
    .B1(_0816_),
    .B2(_0818_),
    .C1(_0819_),
    .X(_0820_));
 sky130_fd_sc_hd__a22o_1 _1377_ (.A1(net67),
    .A2(_0490_),
    .B1(_0491_),
    .B2(net66),
    .X(_0821_));
 sky130_fd_sc_hd__a31o_1 _1378_ (.A1(_0466_),
    .A2(\fast_pwm_inst.pwm_counter[8] ),
    .A3(_0817_),
    .B1(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__or2_1 _1379_ (.A(net66),
    .B(_0491_),
    .X(_0823_));
 sky130_fd_sc_hd__o221a_1 _1380_ (.A1(net67),
    .A2(_0490_),
    .B1(_0820_),
    .B2(_0822_),
    .C1(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _1381_ (.A(_0463_),
    .B(\fast_pwm_inst.pwm_counter[15] ),
    .Y(_0825_));
 sky130_fd_sc_hd__o21ai_1 _1382_ (.A1(net70),
    .A2(_0487_),
    .B1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nor2_1 _1383_ (.A(_0463_),
    .B(\fast_pwm_inst.pwm_counter[15] ),
    .Y(_0827_));
 sky130_fd_sc_hd__a221o_1 _1384_ (.A1(net70),
    .A2(_0487_),
    .B1(_0488_),
    .B2(net69),
    .C1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__or2_1 _1385_ (.A(_0826_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__nor3_1 _1386_ (.A(_0465_),
    .B(\fast_pwm_inst.pwm_counter[11] ),
    .C(_0823_),
    .Y(_0830_));
 sky130_fd_sc_hd__o22a_1 _1387_ (.A1(net69),
    .A2(_0488_),
    .B1(_0489_),
    .B2(net68),
    .X(_0831_));
 sky130_fd_sc_hd__a21o_1 _1388_ (.A1(net68),
    .A2(_0489_),
    .B1(_0824_),
    .X(_0832_));
 sky130_fd_sc_hd__or4b_1 _1389_ (.A(_0829_),
    .B(_0832_),
    .C(_0830_),
    .D_N(_0831_),
    .X(_0833_));
 sky130_fd_sc_hd__o31a_1 _1390_ (.A1(net70),
    .A2(_0487_),
    .A3(_0827_),
    .B1(_0825_),
    .X(_0834_));
 sky130_fd_sc_hd__o211a_1 _1391_ (.A1(_0829_),
    .A2(_0831_),
    .B1(_0833_),
    .C1(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__a21o_1 _1392_ (.A1(net72),
    .A2(_0486_),
    .B1(_0795_),
    .X(_0836_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_0794_),
    .B(_0796_),
    .Y(_0837_));
 sky130_fd_sc_hd__a211o_1 _1394_ (.A1(_0461_),
    .A2(\fast_pwm_inst.pwm_counter[21] ),
    .B1(_0792_),
    .C1(_0793_),
    .X(_0838_));
 sky130_fd_sc_hd__or4b_1 _1395_ (.A(_0836_),
    .B(_0837_),
    .C(_0838_),
    .D_N(_0801_),
    .X(_0839_));
 sky130_fd_sc_hd__o32a_1 _1396_ (.A1(_0800_),
    .A2(_0835_),
    .A3(_0839_),
    .B1(_0804_),
    .B2(_0792_),
    .X(_0840_));
 sky130_fd_sc_hd__o221a_1 _1397_ (.A1(net86),
    .A2(_0473_),
    .B1(_0474_),
    .B2(net85),
    .C1(_0782_),
    .X(_0841_));
 sky130_fd_sc_hd__or3b_1 _1398_ (.A(_0783_),
    .B(_0789_),
    .C_N(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__a21o_1 _1399_ (.A1(net85),
    .A2(_0474_),
    .B1(_0786_),
    .X(_0843_));
 sky130_fd_sc_hd__a211o_1 _1400_ (.A1(net81),
    .A2(_0478_),
    .B1(_0791_),
    .C1(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__o221a_1 _1401_ (.A1(_0458_),
    .A2(\fast_pwm_inst.pwm_counter[25] ),
    .B1(_0478_),
    .B2(net81),
    .C1(_0781_),
    .X(_0845_));
 sky130_fd_sc_hd__or3b_1 _1402_ (.A(_0842_),
    .B(_0844_),
    .C_N(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__o22a_4 _1403_ (.A1(_0790_),
    .A2(_0791_),
    .B1(_0840_),
    .B2(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__and2_1 _1404_ (.A(_0501_),
    .B(_0847_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_1 _1405_ (.A(\fast_pwm_inst.pwm_counter[1] ),
    .B(\fast_pwm_inst.pwm_counter[0] ),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_1 _1406_ (.A(\fast_pwm_inst.pwm_counter[1] ),
    .B(\fast_pwm_inst.pwm_counter[0] ),
    .X(_0849_));
 sky130_fd_sc_hd__and3_1 _1407_ (.A(_0847_),
    .B(_0848_),
    .C(_0849_),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _1408_ (.A(_0499_),
    .B(_0848_),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_1 _1409_ (.A(_0499_),
    .B(_0848_),
    .Y(_0851_));
 sky130_fd_sc_hd__and3b_1 _1410_ (.A_N(_0851_),
    .B(_0847_),
    .C(_0850_),
    .X(_0022_));
 sky130_fd_sc_hd__and4_1 _1411_ (.A(\fast_pwm_inst.pwm_counter[3] ),
    .B(\fast_pwm_inst.pwm_counter[2] ),
    .C(\fast_pwm_inst.pwm_counter[1] ),
    .D(\fast_pwm_inst.pwm_counter[0] ),
    .X(_0852_));
 sky130_fd_sc_hd__or2_1 _1412_ (.A(\fast_pwm_inst.pwm_counter[3] ),
    .B(_0851_),
    .X(_0853_));
 sky130_fd_sc_hd__and3b_1 _1413_ (.A_N(_0852_),
    .B(_0853_),
    .C(_0847_),
    .X(_0025_));
 sky130_fd_sc_hd__nand2_1 _1414_ (.A(\fast_pwm_inst.pwm_counter[4] ),
    .B(_0852_),
    .Y(_0854_));
 sky130_fd_sc_hd__or2_1 _1415_ (.A(\fast_pwm_inst.pwm_counter[4] ),
    .B(_0852_),
    .X(_0855_));
 sky130_fd_sc_hd__and3_1 _1416_ (.A(_0847_),
    .B(_0854_),
    .C(_0855_),
    .X(_0026_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0496_),
    .B(_0854_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _1418_ (.A(_0496_),
    .B(_0854_),
    .Y(_0857_));
 sky130_fd_sc_hd__and3b_1 _1419_ (.A_N(_0856_),
    .B(_0857_),
    .C(_0847_),
    .X(_0027_));
 sky130_fd_sc_hd__and4_1 _1420_ (.A(\fast_pwm_inst.pwm_counter[6] ),
    .B(\fast_pwm_inst.pwm_counter[5] ),
    .C(\fast_pwm_inst.pwm_counter[4] ),
    .D(_0852_),
    .X(_0858_));
 sky130_fd_sc_hd__or2_1 _1421_ (.A(\fast_pwm_inst.pwm_counter[6] ),
    .B(_0856_),
    .X(_0859_));
 sky130_fd_sc_hd__and3b_1 _1422_ (.A_N(_0858_),
    .B(_0859_),
    .C(_0847_),
    .X(_0028_));
 sky130_fd_sc_hd__nand2_1 _1423_ (.A(\fast_pwm_inst.pwm_counter[7] ),
    .B(_0858_),
    .Y(_0860_));
 sky130_fd_sc_hd__or2_1 _1424_ (.A(\fast_pwm_inst.pwm_counter[7] ),
    .B(_0858_),
    .X(_0861_));
 sky130_fd_sc_hd__and3_1 _1425_ (.A(_0847_),
    .B(_0860_),
    .C(_0861_),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _1426_ (.A(_0493_),
    .B(_0860_),
    .Y(_0862_));
 sky130_fd_sc_hd__nand2_1 _1427_ (.A(_0493_),
    .B(_0860_),
    .Y(_0863_));
 sky130_fd_sc_hd__and3b_1 _1428_ (.A_N(_0862_),
    .B(_0863_),
    .C(_0847_),
    .X(_0030_));
 sky130_fd_sc_hd__and4_1 _1429_ (.A(\fast_pwm_inst.pwm_counter[9] ),
    .B(\fast_pwm_inst.pwm_counter[8] ),
    .C(\fast_pwm_inst.pwm_counter[7] ),
    .D(_0858_),
    .X(_0864_));
 sky130_fd_sc_hd__or2_1 _1430_ (.A(\fast_pwm_inst.pwm_counter[9] ),
    .B(_0862_),
    .X(_0865_));
 sky130_fd_sc_hd__and3b_1 _1431_ (.A_N(_0864_),
    .B(_0865_),
    .C(_0847_),
    .X(_0031_));
 sky130_fd_sc_hd__nand2_1 _1432_ (.A(\fast_pwm_inst.pwm_counter[10] ),
    .B(_0864_),
    .Y(_0866_));
 sky130_fd_sc_hd__or2_1 _1433_ (.A(\fast_pwm_inst.pwm_counter[10] ),
    .B(_0864_),
    .X(_0867_));
 sky130_fd_sc_hd__and3_1 _1434_ (.A(_0847_),
    .B(_0866_),
    .C(_0867_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _1435_ (.A(_0490_),
    .B(_0866_),
    .Y(_0868_));
 sky130_fd_sc_hd__nand2_1 _1436_ (.A(_0490_),
    .B(_0866_),
    .Y(_0869_));
 sky130_fd_sc_hd__and3b_1 _1437_ (.A_N(_0868_),
    .B(_0869_),
    .C(_0847_),
    .X(_0002_));
 sky130_fd_sc_hd__and4_1 _1438_ (.A(\fast_pwm_inst.pwm_counter[12] ),
    .B(\fast_pwm_inst.pwm_counter[11] ),
    .C(\fast_pwm_inst.pwm_counter[10] ),
    .D(_0864_),
    .X(_0870_));
 sky130_fd_sc_hd__or2_1 _1439_ (.A(\fast_pwm_inst.pwm_counter[12] ),
    .B(_0868_),
    .X(_0871_));
 sky130_fd_sc_hd__and3b_1 _1440_ (.A_N(_0870_),
    .B(_0871_),
    .C(_0847_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2_1 _1441_ (.A(\fast_pwm_inst.pwm_counter[13] ),
    .B(_0870_),
    .Y(_0872_));
 sky130_fd_sc_hd__or2_1 _1442_ (.A(\fast_pwm_inst.pwm_counter[13] ),
    .B(_0870_),
    .X(_0873_));
 sky130_fd_sc_hd__and3_1 _1443_ (.A(_0847_),
    .B(_0872_),
    .C(_0873_),
    .X(_0004_));
 sky130_fd_sc_hd__nor2_1 _1444_ (.A(_0487_),
    .B(_0872_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_1 _1445_ (.A(_0487_),
    .B(_0872_),
    .Y(_0875_));
 sky130_fd_sc_hd__and3b_1 _1446_ (.A_N(_0874_),
    .B(_0875_),
    .C(_0847_),
    .X(_0005_));
 sky130_fd_sc_hd__and4_1 _1447_ (.A(\fast_pwm_inst.pwm_counter[15] ),
    .B(\fast_pwm_inst.pwm_counter[14] ),
    .C(\fast_pwm_inst.pwm_counter[13] ),
    .D(_0870_),
    .X(_0876_));
 sky130_fd_sc_hd__or2_1 _1448_ (.A(\fast_pwm_inst.pwm_counter[15] ),
    .B(_0874_),
    .X(_0877_));
 sky130_fd_sc_hd__and3b_1 _1449_ (.A_N(_0876_),
    .B(_0877_),
    .C(_0847_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _1450_ (.A(\fast_pwm_inst.pwm_counter[16] ),
    .B(_0876_),
    .Y(_0878_));
 sky130_fd_sc_hd__or2_1 _1451_ (.A(\fast_pwm_inst.pwm_counter[16] ),
    .B(_0876_),
    .X(_0879_));
 sky130_fd_sc_hd__and3_1 _1452_ (.A(_0847_),
    .B(_0878_),
    .C(_0879_),
    .X(_0007_));
 sky130_fd_sc_hd__nor2_1 _1453_ (.A(_0485_),
    .B(_0878_),
    .Y(_0880_));
 sky130_fd_sc_hd__nand2_1 _1454_ (.A(_0485_),
    .B(_0878_),
    .Y(_0881_));
 sky130_fd_sc_hd__and3b_1 _1455_ (.A_N(_0880_),
    .B(_0881_),
    .C(_0847_),
    .X(_0008_));
 sky130_fd_sc_hd__and4_1 _1456_ (.A(\fast_pwm_inst.pwm_counter[18] ),
    .B(\fast_pwm_inst.pwm_counter[17] ),
    .C(\fast_pwm_inst.pwm_counter[16] ),
    .D(_0876_),
    .X(_0882_));
 sky130_fd_sc_hd__or2_1 _1457_ (.A(\fast_pwm_inst.pwm_counter[18] ),
    .B(_0880_),
    .X(_0883_));
 sky130_fd_sc_hd__and3b_1 _1458_ (.A_N(_0882_),
    .B(_0883_),
    .C(_0847_),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(\fast_pwm_inst.pwm_counter[19] ),
    .B(_0882_),
    .Y(_0884_));
 sky130_fd_sc_hd__or2_1 _1460_ (.A(\fast_pwm_inst.pwm_counter[19] ),
    .B(_0882_),
    .X(_0885_));
 sky130_fd_sc_hd__and3_1 _1461_ (.A(_0847_),
    .B(_0884_),
    .C(_0885_),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _1462_ (.A(_0482_),
    .B(_0884_),
    .Y(_0886_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(_0482_),
    .B(_0884_),
    .Y(_0887_));
 sky130_fd_sc_hd__and3b_1 _1464_ (.A_N(_0886_),
    .B(_0887_),
    .C(_0847_),
    .X(_0012_));
 sky130_fd_sc_hd__and4_1 _1465_ (.A(\fast_pwm_inst.pwm_counter[21] ),
    .B(\fast_pwm_inst.pwm_counter[20] ),
    .C(\fast_pwm_inst.pwm_counter[19] ),
    .D(_0882_),
    .X(_0888_));
 sky130_fd_sc_hd__inv_2 _1466_ (.A(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__o211a_1 _1467_ (.A1(\fast_pwm_inst.pwm_counter[21] ),
    .A2(_0886_),
    .B1(_0889_),
    .C1(_0847_),
    .X(_0013_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(\fast_pwm_inst.pwm_counter[22] ),
    .B(_0888_),
    .Y(_0890_));
 sky130_fd_sc_hd__o211a_1 _1469_ (.A1(\fast_pwm_inst.pwm_counter[22] ),
    .A2(_0888_),
    .B1(_0890_),
    .C1(_0847_),
    .X(_0014_));
 sky130_fd_sc_hd__nor2_1 _1470_ (.A(_0479_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _1471_ (.A(_0479_),
    .B(_0890_),
    .Y(_0892_));
 sky130_fd_sc_hd__and3b_1 _1472_ (.A_N(_0891_),
    .B(_0892_),
    .C(_0847_),
    .X(_0015_));
 sky130_fd_sc_hd__and4_1 _1473_ (.A(\fast_pwm_inst.pwm_counter[24] ),
    .B(\fast_pwm_inst.pwm_counter[23] ),
    .C(\fast_pwm_inst.pwm_counter[22] ),
    .D(_0888_),
    .X(_0893_));
 sky130_fd_sc_hd__inv_2 _1474_ (.A(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__o211a_1 _1475_ (.A1(\fast_pwm_inst.pwm_counter[24] ),
    .A2(_0891_),
    .B1(_0894_),
    .C1(_0847_),
    .X(_0016_));
 sky130_fd_sc_hd__or2_1 _1476_ (.A(\fast_pwm_inst.pwm_counter[25] ),
    .B(_0893_),
    .X(_0895_));
 sky130_fd_sc_hd__nor2_1 _1477_ (.A(_0477_),
    .B(_0894_),
    .Y(_0896_));
 sky130_fd_sc_hd__and3b_1 _1478_ (.A_N(_0896_),
    .B(_0847_),
    .C(_0895_),
    .X(_0017_));
 sky130_fd_sc_hd__or2_1 _1479_ (.A(\fast_pwm_inst.pwm_counter[26] ),
    .B(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__and3_1 _1480_ (.A(\fast_pwm_inst.pwm_counter[26] ),
    .B(\fast_pwm_inst.pwm_counter[25] ),
    .C(_0893_),
    .X(_0898_));
 sky130_fd_sc_hd__and3b_1 _1481_ (.A_N(_0898_),
    .B(_0847_),
    .C(_0897_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _1482_ (.A(\fast_pwm_inst.pwm_counter[27] ),
    .B(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__and2_1 _1483_ (.A(\fast_pwm_inst.pwm_counter[27] ),
    .B(_0898_),
    .X(_0900_));
 sky130_fd_sc_hd__and3b_1 _1484_ (.A_N(_0900_),
    .B(_0847_),
    .C(_0899_),
    .X(_0019_));
 sky130_fd_sc_hd__or2_1 _1485_ (.A(\fast_pwm_inst.pwm_counter[28] ),
    .B(_0900_),
    .X(_0901_));
 sky130_fd_sc_hd__nand2_1 _1486_ (.A(\fast_pwm_inst.pwm_counter[28] ),
    .B(_0900_),
    .Y(_0902_));
 sky130_fd_sc_hd__and3_1 _1487_ (.A(_0847_),
    .B(_0901_),
    .C(_0902_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _1488_ (.A(_0473_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__and3_1 _1489_ (.A(\fast_pwm_inst.pwm_counter[29] ),
    .B(\fast_pwm_inst.pwm_counter[28] ),
    .C(_0900_),
    .X(_0904_));
 sky130_fd_sc_hd__and3b_1 _1490_ (.A_N(_0904_),
    .B(_0847_),
    .C(_0903_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _1491_ (.A(\fast_pwm_inst.pwm_counter[30] ),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(\fast_pwm_inst.pwm_counter[30] ),
    .B(_0904_),
    .Y(_0906_));
 sky130_fd_sc_hd__and3_1 _1493_ (.A(_0847_),
    .B(_0905_),
    .C(_0906_),
    .X(_0023_));
 sky130_fd_sc_hd__a21boi_1 _1494_ (.A1(_0471_),
    .A2(_0906_),
    .B1_N(_0847_),
    .Y(_0024_));
 sky130_fd_sc_hd__a21o_1 _1495_ (.A1(_0470_),
    .A2(_0600_),
    .B1(_0615_),
    .X(_0035_));
 sky130_fd_sc_hd__and2b_1 _1496_ (.A_N(net97),
    .B(net98),
    .X(_0907_));
 sky130_fd_sc_hd__and2b_1 _1497_ (.A_N(net98),
    .B(net97),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _1498_ (.A1(\phase_pwm_inst.pwm_outb ),
    .A2(_0907_),
    .B1(_0908_),
    .B2(\fast_pwm_inst.pwm_outb ),
    .X(net101));
 sky130_fd_sc_hd__a22o_2 _1499_ (.A1(\phase_pwm_inst.pwm_outa ),
    .A2(_0907_),
    .B1(_0908_),
    .B2(\fast_pwm_inst.pwm_outa ),
    .X(net100));
 sky130_fd_sc_hd__a22o_1 _1500_ (.A1(\fast_pwm_inst.pwm_counter[23] ),
    .A2(_0505_),
    .B1(_0506_),
    .B2(\fast_pwm_inst.pwm_counter[22] ),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _1501_ (.A1(_0480_),
    .A2(net47),
    .B1(net46),
    .B2(_0481_),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _1502_ (.A1(\fast_pwm_inst.pwm_counter[19] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(\fast_pwm_inst.pwm_counter[18] ),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _1503_ (.A1(\fast_pwm_inst.pwm_counter[17] ),
    .A2(_0511_),
    .B1(_0512_),
    .B2(\fast_pwm_inst.pwm_counter[16] ),
    .C1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__o22a_1 _1504_ (.A1(\fast_pwm_inst.pwm_counter[20] ),
    .A2(_0508_),
    .B1(_0509_),
    .B2(\fast_pwm_inst.pwm_counter[19] ),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _1505_ (.A1(_0484_),
    .A2(net42),
    .B1(net41),
    .B2(_0485_),
    .X(_0914_));
 sky130_fd_sc_hd__and3b_1 _1506_ (.A_N(_0914_),
    .B(_0912_),
    .C(_0913_),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _1507_ (.A1(\fast_pwm_inst.pwm_counter[21] ),
    .A2(_0507_),
    .B1(_0508_),
    .B2(\fast_pwm_inst.pwm_counter[20] ),
    .X(_0916_));
 sky130_fd_sc_hd__a21o_1 _1508_ (.A1(_0911_),
    .A2(_0913_),
    .B1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__o21ba_1 _1509_ (.A1(_0915_),
    .A2(_0917_),
    .B1_N(_0910_),
    .X(_0918_));
 sky130_fd_sc_hd__a2bb2o_1 _1510_ (.A1_N(_0909_),
    .A2_N(_0918_),
    .B1(_0479_),
    .B2(net48),
    .X(_0919_));
 sky130_fd_sc_hd__nand2_1 _1511_ (.A(\fast_pwm_inst.pwm_counter[3] ),
    .B(_0519_),
    .Y(_0920_));
 sky130_fd_sc_hd__a22o_1 _1512_ (.A1(_0500_),
    .A2(net44),
    .B1(net33),
    .B2(_0501_),
    .X(_0921_));
 sky130_fd_sc_hd__o22a_1 _1513_ (.A1(_0499_),
    .A2(net55),
    .B1(net44),
    .B2(_0500_),
    .X(_0922_));
 sky130_fd_sc_hd__a22o_1 _1514_ (.A1(_0499_),
    .A2(net55),
    .B1(_0921_),
    .B2(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_1 _1515_ (.A(\fast_pwm_inst.pwm_counter[3] ),
    .B(_0519_),
    .Y(_0924_));
 sky130_fd_sc_hd__a221o_1 _1516_ (.A1(_0497_),
    .A2(net59),
    .B1(_0920_),
    .B2(_0923_),
    .C1(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__o22a_1 _1517_ (.A1(_0496_),
    .A2(net60),
    .B1(net59),
    .B2(_0497_),
    .X(_0926_));
 sky130_fd_sc_hd__a22o_1 _1518_ (.A1(_0495_),
    .A2(net61),
    .B1(net60),
    .B2(_0496_),
    .X(_0927_));
 sky130_fd_sc_hd__a21o_1 _1519_ (.A1(_0925_),
    .A2(_0926_),
    .B1(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__o22a_1 _1520_ (.A1(_0494_),
    .A2(net62),
    .B1(net61),
    .B2(_0495_),
    .X(_0929_));
 sky130_fd_sc_hd__a22o_1 _1521_ (.A1(_0493_),
    .A2(net63),
    .B1(net62),
    .B2(_0494_),
    .X(_0930_));
 sky130_fd_sc_hd__a21o_1 _1522_ (.A1(_0928_),
    .A2(_0929_),
    .B1(_0930_),
    .X(_0931_));
 sky130_fd_sc_hd__o221a_1 _1523_ (.A1(_0492_),
    .A2(net64),
    .B1(net63),
    .B2(_0493_),
    .C1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__nor2_1 _1524_ (.A(\fast_pwm_inst.pwm_counter[10] ),
    .B(_0518_),
    .Y(_0933_));
 sky130_fd_sc_hd__a221o_1 _1525_ (.A1(_0490_),
    .A2(net35),
    .B1(net64),
    .B2(_0492_),
    .C1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__nand2_1 _1526_ (.A(\fast_pwm_inst.pwm_counter[10] ),
    .B(_0518_),
    .Y(_0935_));
 sky130_fd_sc_hd__o221a_1 _1527_ (.A1(_0490_),
    .A2(net35),
    .B1(_0932_),
    .B2(_0934_),
    .C1(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__and2_1 _1528_ (.A(\fast_pwm_inst.pwm_counter[15] ),
    .B(_0513_),
    .X(_0937_));
 sky130_fd_sc_hd__nor2_1 _1529_ (.A(\fast_pwm_inst.pwm_counter[15] ),
    .B(_0513_),
    .Y(_0938_));
 sky130_fd_sc_hd__a22o_1 _1530_ (.A1(\fast_pwm_inst.pwm_counter[13] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(\fast_pwm_inst.pwm_counter[12] ),
    .X(_0939_));
 sky130_fd_sc_hd__a221o_1 _1531_ (.A1(_0487_),
    .A2(net38),
    .B1(net37),
    .B2(_0488_),
    .C1(_0938_),
    .X(_0940_));
 sky130_fd_sc_hd__a211o_1 _1532_ (.A1(\fast_pwm_inst.pwm_counter[14] ),
    .A2(_0514_),
    .B1(_0937_),
    .C1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o32ai_1 _1533_ (.A1(\fast_pwm_inst.pwm_counter[11] ),
    .A2(_0517_),
    .A3(_0935_),
    .B1(_0516_),
    .B2(\fast_pwm_inst.pwm_counter[12] ),
    .Y(_0204_));
 sky130_fd_sc_hd__or4_1 _1534_ (.A(_0936_),
    .B(_0939_),
    .C(_0941_),
    .D(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__nand2b_1 _1535_ (.A_N(_0941_),
    .B(_0939_),
    .Y(_0206_));
 sky130_fd_sc_hd__or3_1 _1536_ (.A(_0487_),
    .B(net38),
    .C(_0938_),
    .X(_0207_));
 sky130_fd_sc_hd__and4b_1 _1537_ (.A_N(_0937_),
    .B(_0205_),
    .C(_0206_),
    .D(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a221o_1 _1538_ (.A1(_0479_),
    .A2(net48),
    .B1(net40),
    .B2(_0486_),
    .C1(_0909_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _1539_ (.A(_0914_),
    .B(_0916_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand3b_1 _1540_ (.A_N(_0910_),
    .B(_0913_),
    .C(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__or4_1 _1541_ (.A(_0912_),
    .B(_0208_),
    .C(_0209_),
    .D(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__a2bb2o_1 _1542_ (.A1_N(_0474_),
    .A2_N(net53),
    .B1(_0502_),
    .B2(\fast_pwm_inst.pwm_counter[27] ),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _1543_ (.A1(_0475_),
    .A2(net52),
    .B1(net51),
    .B2(_0476_),
    .X(_0214_));
 sky130_fd_sc_hd__o22a_1 _1544_ (.A1(_0472_),
    .A2(net56),
    .B1(net54),
    .B2(_0473_),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _1545_ (.A1(\fast_pwm_inst.pwm_counter[25] ),
    .A2(_0503_),
    .B1(_0504_),
    .B2(\fast_pwm_inst.pwm_counter[24] ),
    .X(_0216_));
 sky130_fd_sc_hd__or3b_1 _1546_ (.A(_0213_),
    .B(_0214_),
    .C_N(_0215_),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _1547_ (.A1(_0471_),
    .A2(net57),
    .B1(net56),
    .B2(_0472_),
    .X(_0218_));
 sky130_fd_sc_hd__a221o_1 _1548_ (.A1(_0473_),
    .A2(net54),
    .B1(net53),
    .B2(_0474_),
    .C1(_0218_),
    .X(_0219_));
 sky130_fd_sc_hd__or2_1 _1549_ (.A(_0476_),
    .B(net51),
    .X(_0220_));
 sky130_fd_sc_hd__o21ai_1 _1550_ (.A1(\fast_pwm_inst.pwm_counter[24] ),
    .A2(_0504_),
    .B1(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__or4_1 _1551_ (.A(_0216_),
    .B(_0217_),
    .C(_0219_),
    .D(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__a221o_1 _1552_ (.A1(_0477_),
    .A2(net50),
    .B1(_0919_),
    .B2(_0212_),
    .C1(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__o21ai_1 _1553_ (.A1(\fast_pwm_inst.pwm_counter[25] ),
    .A2(_0503_),
    .B1(_0216_),
    .Y(_0224_));
 sky130_fd_sc_hd__a21oi_1 _1554_ (.A1(_0220_),
    .A2(_0224_),
    .B1(_0214_),
    .Y(_0225_));
 sky130_fd_sc_hd__nor2_1 _1555_ (.A(_0213_),
    .B(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__o22a_1 _1556_ (.A1(_0471_),
    .A2(net57),
    .B1(_0219_),
    .B2(_0226_),
    .X(_0227_));
 sky130_fd_sc_hd__o211a_1 _1557_ (.A1(_0215_),
    .A2(_0218_),
    .B1(_0223_),
    .C1(_0227_),
    .X(_0033_));
 sky130_fd_sc_hd__nor2_1 _1558_ (.A(\fast_pwm_inst.pwm_counter[15] ),
    .B(_0532_),
    .Y(_0228_));
 sky130_fd_sc_hd__a22o_1 _1559_ (.A1(\fast_pwm_inst.pwm_counter[15] ),
    .A2(_0532_),
    .B1(_0533_),
    .B2(\fast_pwm_inst.pwm_counter[14] ),
    .X(_0229_));
 sky130_fd_sc_hd__o22a_1 _1560_ (.A1(\fast_pwm_inst.pwm_counter[14] ),
    .A2(_0533_),
    .B1(_0534_),
    .B2(\fast_pwm_inst.pwm_counter[13] ),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _1561_ (.A1(_0487_),
    .A2(net6),
    .B1(net5),
    .B2(_0488_),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _1562_ (.A1(\fast_pwm_inst.pwm_counter[13] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\fast_pwm_inst.pwm_counter[12] ),
    .X(_0232_));
 sky130_fd_sc_hd__a21oi_1 _1563_ (.A1(_0230_),
    .A2(_0232_),
    .B1(_0229_),
    .Y(_0233_));
 sky130_fd_sc_hd__and2_1 _1564_ (.A(_0499_),
    .B(net23),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _1565_ (.A1(_0500_),
    .A2(net12),
    .B1(net1),
    .B2(_0501_),
    .X(_0235_));
 sky130_fd_sc_hd__o221a_1 _1566_ (.A1(_0499_),
    .A2(net23),
    .B1(net12),
    .B2(_0500_),
    .C1(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__o22a_1 _1567_ (.A1(_0498_),
    .A2(net26),
    .B1(_0234_),
    .B2(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__a221o_1 _1568_ (.A1(_0497_),
    .A2(net27),
    .B1(net26),
    .B2(_0498_),
    .C1(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _1569_ (.A1(_0495_),
    .A2(net29),
    .B1(net28),
    .B2(_0496_),
    .X(_0239_));
 sky130_fd_sc_hd__o22a_1 _1570_ (.A1(_0496_),
    .A2(net28),
    .B1(net27),
    .B2(_0497_),
    .X(_0240_));
 sky130_fd_sc_hd__a21o_1 _1571_ (.A1(_0238_),
    .A2(_0240_),
    .B1(_0239_),
    .X(_0241_));
 sky130_fd_sc_hd__o22a_1 _1572_ (.A1(_0494_),
    .A2(net30),
    .B1(net29),
    .B2(_0495_),
    .X(_0242_));
 sky130_fd_sc_hd__a22o_1 _1573_ (.A1(_0493_),
    .A2(net31),
    .B1(net30),
    .B2(_0494_),
    .X(_0243_));
 sky130_fd_sc_hd__a21o_1 _1574_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o22a_1 _1575_ (.A1(_0492_),
    .A2(net32),
    .B1(net31),
    .B2(_0493_),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _1576_ (.A1(_0491_),
    .A2(net2),
    .B1(net32),
    .B2(_0492_),
    .X(_0246_));
 sky130_fd_sc_hd__a21o_1 _1577_ (.A1(_0244_),
    .A2(_0245_),
    .B1(_0246_),
    .X(_0247_));
 sky130_fd_sc_hd__o221a_1 _1578_ (.A1(_0490_),
    .A2(net3),
    .B1(net2),
    .B2(_0491_),
    .C1(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__a221o_1 _1579_ (.A1(_0489_),
    .A2(net4),
    .B1(net3),
    .B2(_0490_),
    .C1(_0228_),
    .X(_0249_));
 sky130_fd_sc_hd__or4_1 _1580_ (.A(_0229_),
    .B(_0231_),
    .C(_0232_),
    .D(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__o22a_1 _1581_ (.A1(_0228_),
    .A2(_0233_),
    .B1(_0248_),
    .B2(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _1582_ (.A1(_0480_),
    .A2(net15),
    .B1(net14),
    .B2(_0481_),
    .X(_0252_));
 sky130_fd_sc_hd__a22o_1 _1583_ (.A1(_0483_),
    .A2(net11),
    .B1(net10),
    .B2(_0484_),
    .X(_0253_));
 sky130_fd_sc_hd__nor2_1 _1584_ (.A(\fast_pwm_inst.pwm_counter[20] ),
    .B(_0527_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _1585_ (.A(_0485_),
    .B(net9),
    .Y(_0255_));
 sky130_fd_sc_hd__a22o_1 _1586_ (.A1(\fast_pwm_inst.pwm_counter[17] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\fast_pwm_inst.pwm_counter[16] ),
    .X(_0256_));
 sky130_fd_sc_hd__a221o_1 _1587_ (.A1(\fast_pwm_inst.pwm_counter[21] ),
    .A2(_0526_),
    .B1(net8),
    .B2(_0486_),
    .C1(_0254_),
    .X(_0257_));
 sky130_fd_sc_hd__a221o_1 _1588_ (.A1(\fast_pwm_inst.pwm_counter[20] ),
    .A2(_0527_),
    .B1(_0528_),
    .B2(\fast_pwm_inst.pwm_counter[19] ),
    .C1(_0253_),
    .X(_0258_));
 sky130_fd_sc_hd__or4_1 _1589_ (.A(_0252_),
    .B(_0256_),
    .C(_0257_),
    .D(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__a221o_1 _1590_ (.A1(\fast_pwm_inst.pwm_counter[18] ),
    .A2(_0529_),
    .B1(net9),
    .B2(_0485_),
    .C1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__o22a_1 _1591_ (.A1(_0479_),
    .A2(net16),
    .B1(net15),
    .B2(_0480_),
    .X(_0261_));
 sky130_fd_sc_hd__o2bb2a_1 _1592_ (.A1_N(_0255_),
    .A2_N(_0256_),
    .B1(_0484_),
    .B2(net10),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _1593_ (.A(_0253_),
    .B(_0262_),
    .X(_0263_));
 sky130_fd_sc_hd__o221a_1 _1594_ (.A1(_0482_),
    .A2(net13),
    .B1(net11),
    .B2(_0483_),
    .C1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__o22a_1 _1595_ (.A1(_0481_),
    .A2(net14),
    .B1(_0254_),
    .B2(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _1596_ (.A(_0252_),
    .B(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o211a_1 _1597_ (.A1(_0251_),
    .A2(_0260_),
    .B1(_0261_),
    .C1(_0266_),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _1598_ (.A1(_0471_),
    .A2(net25),
    .B1(net24),
    .B2(_0472_),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _1599_ (.A1(\fast_pwm_inst.pwm_counter[28] ),
    .A2(_0521_),
    .B1(_0522_),
    .B2(\fast_pwm_inst.pwm_counter[27] ),
    .X(_0269_));
 sky130_fd_sc_hd__o22a_1 _1600_ (.A1(_0472_),
    .A2(net24),
    .B1(net22),
    .B2(_0473_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _1601_ (.A1(\fast_pwm_inst.pwm_counter[25] ),
    .A2(_0524_),
    .B1(_0525_),
    .B2(\fast_pwm_inst.pwm_counter[24] ),
    .X(_0271_));
 sky130_fd_sc_hd__or3b_1 _1602_ (.A(_0268_),
    .B(_0269_),
    .C_N(_0270_),
    .X(_0272_));
 sky130_fd_sc_hd__o22a_1 _1603_ (.A1(\fast_pwm_inst.pwm_counter[29] ),
    .A2(_0520_),
    .B1(_0521_),
    .B2(\fast_pwm_inst.pwm_counter[28] ),
    .X(_0273_));
 sky130_fd_sc_hd__o221a_1 _1604_ (.A1(\fast_pwm_inst.pwm_counter[27] ),
    .A2(_0522_),
    .B1(_0523_),
    .B2(\fast_pwm_inst.pwm_counter[26] ),
    .C1(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__o2bb2a_1 _1605_ (.A1_N(net16),
    .A2_N(_0479_),
    .B1(\fast_pwm_inst.pwm_counter[24] ),
    .B2(_0525_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_1 _1606_ (.A(_0477_),
    .B(net18),
    .Y(_0276_));
 sky130_fd_sc_hd__o2111a_1 _1607_ (.A1(_0476_),
    .A2(net19),
    .B1(_0274_),
    .C1(_0275_),
    .D1(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__or4b_1 _1608_ (.A(_0267_),
    .B(_0271_),
    .C(_0272_),
    .D_N(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__a22o_1 _1609_ (.A1(\fast_pwm_inst.pwm_counter[26] ),
    .A2(_0523_),
    .B1(_0271_),
    .B2(_0276_),
    .X(_0279_));
 sky130_fd_sc_hd__a21bo_1 _1610_ (.A1(_0269_),
    .A2(_0273_),
    .B1_N(_0270_),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_1 _1611_ (.A1(_0274_),
    .A2(_0279_),
    .B1(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__o221a_1 _1612_ (.A1(_0471_),
    .A2(net25),
    .B1(_0268_),
    .B2(_0281_),
    .C1(_0278_),
    .X(_0032_));
 sky130_fd_sc_hd__a22o_1 _1613_ (.A1(\phase_pwm_inst.counter[13] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(\phase_pwm_inst.counter[12] ),
    .X(_0282_));
 sky130_fd_sc_hd__o21ai_1 _1614_ (.A1(\phase_pwm_inst.counter[13] ),
    .A2(_0515_),
    .B1(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__or2_1 _1615_ (.A(_0446_),
    .B(net60),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _1616_ (.A1(_0450_),
    .A2(net44),
    .B1(net33),
    .B2(_0451_),
    .X(_0285_));
 sky130_fd_sc_hd__o22a_1 _1617_ (.A1(_0449_),
    .A2(net55),
    .B1(net44),
    .B2(_0450_),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _1618_ (.A1(_0448_),
    .A2(net58),
    .B1(net55),
    .B2(_0449_),
    .X(_0287_));
 sky130_fd_sc_hd__a21o_1 _1619_ (.A1(_0285_),
    .A2(_0286_),
    .B1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__o22a_1 _1620_ (.A1(_0447_),
    .A2(net59),
    .B1(net58),
    .B2(_0448_),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _1621_ (.A1(_0446_),
    .A2(net60),
    .B1(net59),
    .B2(_0447_),
    .X(_0290_));
 sky130_fd_sc_hd__a21o_1 _1622_ (.A1(_0288_),
    .A2(_0289_),
    .B1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _1623_ (.A1(_0445_),
    .A2(net61),
    .B1(_0284_),
    .B2(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__o22a_1 _1624_ (.A1(_0444_),
    .A2(net62),
    .B1(net61),
    .B2(_0445_),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _1625_ (.A1(_0443_),
    .A2(net63),
    .B1(net62),
    .B2(_0444_),
    .X(_0294_));
 sky130_fd_sc_hd__a21o_1 _1626_ (.A1(_0292_),
    .A2(_0293_),
    .B1(_0294_),
    .X(_0295_));
 sky130_fd_sc_hd__o22a_1 _1627_ (.A1(_0442_),
    .A2(net64),
    .B1(net63),
    .B2(_0443_),
    .X(_0296_));
 sky130_fd_sc_hd__a22o_1 _1628_ (.A1(_0441_),
    .A2(net34),
    .B1(net64),
    .B2(_0442_),
    .X(_0297_));
 sky130_fd_sc_hd__a21o_1 _1629_ (.A1(_0295_),
    .A2(_0296_),
    .B1(_0297_),
    .X(_0298_));
 sky130_fd_sc_hd__o22a_1 _1630_ (.A1(_0440_),
    .A2(net35),
    .B1(net34),
    .B2(_0441_),
    .X(_0299_));
 sky130_fd_sc_hd__o22a_1 _1631_ (.A1(\phase_pwm_inst.counter[13] ),
    .A2(_0515_),
    .B1(_0516_),
    .B2(\phase_pwm_inst.counter[12] ),
    .X(_0300_));
 sky130_fd_sc_hd__o21ai_1 _1632_ (.A1(\phase_pwm_inst.counter[11] ),
    .A2(_0517_),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__a211o_1 _1633_ (.A1(_0298_),
    .A2(_0299_),
    .B1(_0301_),
    .C1(_0282_),
    .X(_0302_));
 sky130_fd_sc_hd__a22o_1 _1634_ (.A1(_0438_),
    .A2(net38),
    .B1(_0283_),
    .B2(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__o221ai_2 _1635_ (.A1(_0437_),
    .A2(net39),
    .B1(net38),
    .B2(_0438_),
    .C1(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__a22o_1 _1636_ (.A1(\phase_pwm_inst.counter[21] ),
    .A2(_0507_),
    .B1(_0508_),
    .B2(\phase_pwm_inst.counter[20] ),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _1637_ (.A1(_0432_),
    .A2(net45),
    .B1(net43),
    .B2(_0433_),
    .C1(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_1 _1638_ (.A1(_0434_),
    .A2(net42),
    .B1(net41),
    .B2(_0435_),
    .C1(_0306_),
    .X(_0307_));
 sky130_fd_sc_hd__nor2_1 _1639_ (.A(\phase_pwm_inst.counter[23] ),
    .B(_0505_),
    .Y(_0308_));
 sky130_fd_sc_hd__a221o_1 _1640_ (.A1(_0430_),
    .A2(net47),
    .B1(net46),
    .B2(_0431_),
    .C1(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _1641_ (.A1(\phase_pwm_inst.counter[19] ),
    .A2(_0509_),
    .B1(_0510_),
    .B2(\phase_pwm_inst.counter[18] ),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _1642_ (.A1(\phase_pwm_inst.counter[17] ),
    .A2(_0511_),
    .B1(_0512_),
    .B2(\phase_pwm_inst.counter[16] ),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _1643_ (.A1(\phase_pwm_inst.counter[23] ),
    .A2(_0505_),
    .B1(_0506_),
    .B2(\phase_pwm_inst.counter[22] ),
    .X(_0312_));
 sky130_fd_sc_hd__a221o_1 _1644_ (.A1(_0436_),
    .A2(net40),
    .B1(net39),
    .B2(_0437_),
    .C1(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__or3_1 _1645_ (.A(_0310_),
    .B(_0311_),
    .C(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__nor3_1 _1646_ (.A(_0307_),
    .B(_0309_),
    .C(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2b_1 _1647_ (.A_N(_0308_),
    .B(_0312_),
    .Y(_0316_));
 sky130_fd_sc_hd__o221a_1 _1648_ (.A1(\phase_pwm_inst.counter[18] ),
    .A2(_0510_),
    .B1(_0511_),
    .B2(\phase_pwm_inst.counter[17] ),
    .C1(_0311_),
    .X(_0317_));
 sky130_fd_sc_hd__or2_1 _1649_ (.A(_0310_),
    .B(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__o221a_1 _1650_ (.A1(\phase_pwm_inst.counter[20] ),
    .A2(_0508_),
    .B1(_0509_),
    .B2(\phase_pwm_inst.counter[19] ),
    .C1(_0318_),
    .X(_0319_));
 sky130_fd_sc_hd__nor2_1 _1651_ (.A(_0305_),
    .B(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_1 _1652_ (.A1(_0309_),
    .A2(_0320_),
    .B1(_0316_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21oi_1 _1653_ (.A1(_0304_),
    .A2(_0315_),
    .B1(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__a22o_1 _1654_ (.A1(_0423_),
    .A2(net54),
    .B1(net53),
    .B2(_0424_),
    .X(_0323_));
 sky130_fd_sc_hd__a22o_1 _1655_ (.A1(\phase_pwm_inst.counter[25] ),
    .A2(_0503_),
    .B1(_0504_),
    .B2(\phase_pwm_inst.counter[24] ),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _1656_ (.A1(_0421_),
    .A2(net57),
    .B1(net56),
    .B2(_0422_),
    .X(_0325_));
 sky130_fd_sc_hd__o22ai_1 _1657_ (.A1(_0422_),
    .A2(net56),
    .B1(net54),
    .B2(_0423_),
    .Y(_0326_));
 sky130_fd_sc_hd__or4_1 _1658_ (.A(_0323_),
    .B(_0324_),
    .C(_0325_),
    .D(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__o22a_1 _1659_ (.A1(_0425_),
    .A2(net52),
    .B1(net51),
    .B2(_0426_),
    .X(_0328_));
 sky130_fd_sc_hd__nor2_1 _1660_ (.A(\phase_pwm_inst.counter[27] ),
    .B(_0502_),
    .Y(_0329_));
 sky130_fd_sc_hd__a21oi_1 _1661_ (.A1(_0426_),
    .A2(net51),
    .B1(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _1662_ (.A(_0328_),
    .B(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_1 _1663_ (.A(_0424_),
    .B(net53),
    .Y(_0332_));
 sky130_fd_sc_hd__a221o_1 _1664_ (.A1(_0427_),
    .A2(net50),
    .B1(net49),
    .B2(_0428_),
    .C1(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__or4_1 _1665_ (.A(_0322_),
    .B(_0327_),
    .C(_0331_),
    .D(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__o21ai_1 _1666_ (.A1(\phase_pwm_inst.counter[25] ),
    .A2(_0503_),
    .B1(_0324_),
    .Y(_0335_));
 sky130_fd_sc_hd__or2_1 _1667_ (.A(_0328_),
    .B(_0329_),
    .X(_0336_));
 sky130_fd_sc_hd__o221a_1 _1668_ (.A1(_0424_),
    .A2(net53),
    .B1(_0331_),
    .B2(_0335_),
    .C1(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o21ba_1 _1669_ (.A1(_0323_),
    .A2(_0337_),
    .B1_N(_0326_),
    .X(_0338_));
 sky130_fd_sc_hd__o221a_1 _1670_ (.A1(_0421_),
    .A2(net57),
    .B1(_0325_),
    .B2(_0338_),
    .C1(_0334_),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _1671_ (.A1(_0421_),
    .A2(net25),
    .B1(net24),
    .B2(_0422_),
    .X(_0339_));
 sky130_fd_sc_hd__a2bb2o_1 _1672_ (.A1_N(_0422_),
    .A2_N(net24),
    .B1(_0520_),
    .B2(\phase_pwm_inst.counter[29] ),
    .X(_0340_));
 sky130_fd_sc_hd__o22a_1 _1673_ (.A1(\phase_pwm_inst.counter[29] ),
    .A2(_0520_),
    .B1(_0521_),
    .B2(\phase_pwm_inst.counter[28] ),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _1674_ (.A1(\phase_pwm_inst.counter[28] ),
    .A2(_0521_),
    .B1(_0522_),
    .B2(\phase_pwm_inst.counter[27] ),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _1675_ (.A1(\phase_pwm_inst.counter[26] ),
    .A2(_0523_),
    .B1(_0524_),
    .B2(\phase_pwm_inst.counter[25] ),
    .X(_0343_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(_0427_),
    .B(net18),
    .Y(_0344_));
 sky130_fd_sc_hd__a31o_1 _1677_ (.A1(\phase_pwm_inst.counter[24] ),
    .A2(_0525_),
    .A3(_0344_),
    .B1(_0343_),
    .X(_0345_));
 sky130_fd_sc_hd__o221a_1 _1678_ (.A1(\phase_pwm_inst.counter[27] ),
    .A2(_0522_),
    .B1(_0523_),
    .B2(\phase_pwm_inst.counter[26] ),
    .C1(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__or2_1 _1679_ (.A(_0342_),
    .B(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__a21oi_1 _1680_ (.A1(_0341_),
    .A2(_0347_),
    .B1(_0340_),
    .Y(_0348_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(_0429_),
    .A2(net16),
    .B1(net15),
    .B2(_0430_),
    .X(_0349_));
 sky130_fd_sc_hd__o21a_1 _1682_ (.A1(_0429_),
    .A2(net16),
    .B1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _1683_ (.A1(_0431_),
    .A2(net14),
    .B1(net13),
    .B2(_0432_),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_1 _1684_ (.A1(\phase_pwm_inst.counter[17] ),
    .A2(_0530_),
    .B1(_0531_),
    .B2(\phase_pwm_inst.counter[16] ),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _1685_ (.A1(\phase_pwm_inst.counter[19] ),
    .A2(_0528_),
    .B1(_0529_),
    .B2(\phase_pwm_inst.counter[18] ),
    .X(_0353_));
 sky130_fd_sc_hd__inv_2 _1686_ (.A(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(\phase_pwm_inst.counter[19] ),
    .B(_0528_),
    .Y(_0355_));
 sky130_fd_sc_hd__a221o_1 _1688_ (.A1(_0434_),
    .A2(net10),
    .B1(net9),
    .B2(_0435_),
    .C1(_0355_),
    .X(_0356_));
 sky130_fd_sc_hd__or3b_1 _1689_ (.A(_0353_),
    .B(_0356_),
    .C_N(_0352_),
    .X(_0357_));
 sky130_fd_sc_hd__o221a_1 _1690_ (.A1(_0432_),
    .A2(net13),
    .B1(_0354_),
    .B2(_0355_),
    .C1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__o22a_1 _1691_ (.A1(_0429_),
    .A2(net16),
    .B1(net14),
    .B2(_0431_),
    .X(_0359_));
 sky130_fd_sc_hd__nor2_1 _1692_ (.A(_0430_),
    .B(net15),
    .Y(_0360_));
 sky130_fd_sc_hd__o221a_1 _1693_ (.A1(_0430_),
    .A2(net15),
    .B1(_0351_),
    .B2(_0358_),
    .C1(_0359_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2b_1 _1694_ (.A_N(net26),
    .B(\phase_pwm_inst.counter[3] ),
    .Y(_0362_));
 sky130_fd_sc_hd__a22o_1 _1695_ (.A1(_0450_),
    .A2(net12),
    .B1(net1),
    .B2(_0451_),
    .X(_0363_));
 sky130_fd_sc_hd__o22a_1 _1696_ (.A1(_0449_),
    .A2(net23),
    .B1(net12),
    .B2(_0450_),
    .X(_0364_));
 sky130_fd_sc_hd__and2b_1 _1697_ (.A_N(\phase_pwm_inst.counter[3] ),
    .B(net26),
    .X(_0365_));
 sky130_fd_sc_hd__a221o_1 _1698_ (.A1(_0449_),
    .A2(net23),
    .B1(_0363_),
    .B2(_0364_),
    .C1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__a22o_1 _1699_ (.A1(_0447_),
    .A2(net27),
    .B1(_0362_),
    .B2(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_1 _1700_ (.A1(_0446_),
    .A2(net28),
    .B1(net27),
    .B2(_0447_),
    .X(_0368_));
 sky130_fd_sc_hd__a22o_1 _1701_ (.A1(_0445_),
    .A2(net29),
    .B1(net28),
    .B2(_0446_),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _1702_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__o221a_1 _1703_ (.A1(_0444_),
    .A2(net30),
    .B1(net29),
    .B2(_0445_),
    .C1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _1704_ (.A1(_0443_),
    .A2(net31),
    .B1(net30),
    .B2(_0444_),
    .X(_0372_));
 sky130_fd_sc_hd__o22a_1 _1705_ (.A1(_0442_),
    .A2(net32),
    .B1(net31),
    .B2(_0443_),
    .X(_0373_));
 sky130_fd_sc_hd__o21a_1 _1706_ (.A1(_0371_),
    .A2(_0372_),
    .B1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _1707_ (.A1(_0441_),
    .A2(net2),
    .B1(net32),
    .B2(_0442_),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _1708_ (.A(_0440_),
    .B(net3),
    .X(_0376_));
 sky130_fd_sc_hd__a211o_1 _1709_ (.A1(\phase_pwm_inst.counter[10] ),
    .A2(_0536_),
    .B1(_0375_),
    .C1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__or2_1 _1710_ (.A(net2),
    .B(_0376_),
    .X(_0378_));
 sky130_fd_sc_hd__o22a_1 _1711_ (.A1(_0440_),
    .A2(net3),
    .B1(_0378_),
    .B2(_0441_),
    .X(_0379_));
 sky130_fd_sc_hd__o21a_1 _1712_ (.A1(_0374_),
    .A2(_0377_),
    .B1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__nor2_1 _1713_ (.A(_0437_),
    .B(net7),
    .Y(_0381_));
 sky130_fd_sc_hd__a21o_1 _1714_ (.A1(\phase_pwm_inst.counter[14] ),
    .A2(_0533_),
    .B1(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nor2_1 _1715_ (.A(\phase_pwm_inst.counter[15] ),
    .B(_0532_),
    .Y(_0383_));
 sky130_fd_sc_hd__a211o_1 _1716_ (.A1(_0438_),
    .A2(net6),
    .B1(_0382_),
    .C1(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(\phase_pwm_inst.counter[13] ),
    .A2(_0534_),
    .B1(_0535_),
    .B2(\phase_pwm_inst.counter[12] ),
    .X(_0385_));
 sky130_fd_sc_hd__nor2_1 _1718_ (.A(\phase_pwm_inst.counter[13] ),
    .B(_0534_),
    .Y(_0386_));
 sky130_fd_sc_hd__a211o_1 _1719_ (.A1(_0439_),
    .A2(net4),
    .B1(_0385_),
    .C1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__or3_1 _1720_ (.A(_0380_),
    .B(_0384_),
    .C(_0387_),
    .X(_0388_));
 sky130_fd_sc_hd__or3b_1 _1721_ (.A(_0386_),
    .B(_0384_),
    .C_N(_0385_),
    .X(_0389_));
 sky130_fd_sc_hd__or3b_1 _1722_ (.A(net6),
    .B(_0383_),
    .C_N(\phase_pwm_inst.counter[14] ),
    .X(_0390_));
 sky130_fd_sc_hd__and4b_1 _1723_ (.A_N(_0381_),
    .B(_0388_),
    .C(_0389_),
    .D(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__or4b_1 _1724_ (.A(_0349_),
    .B(_0351_),
    .C(_0352_),
    .D_N(_0359_),
    .X(_0392_));
 sky130_fd_sc_hd__a221o_1 _1725_ (.A1(\phase_pwm_inst.counter[20] ),
    .A2(_0527_),
    .B1(net8),
    .B2(_0436_),
    .C1(_0360_),
    .X(_0393_));
 sky130_fd_sc_hd__or4_1 _1726_ (.A(_0353_),
    .B(_0356_),
    .C(_0392_),
    .D(_0393_),
    .X(_0394_));
 sky130_fd_sc_hd__o22a_1 _1727_ (.A1(_0350_),
    .A2(_0361_),
    .B1(_0391_),
    .B2(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__a221o_1 _1728_ (.A1(_0427_),
    .A2(net18),
    .B1(net17),
    .B2(_0428_),
    .C1(_0340_),
    .X(_0396_));
 sky130_fd_sc_hd__a221o_1 _1729_ (.A1(_0425_),
    .A2(net20),
    .B1(net19),
    .B2(_0426_),
    .C1(_0342_),
    .X(_0397_));
 sky130_fd_sc_hd__a221o_1 _1730_ (.A1(_0423_),
    .A2(net22),
    .B1(net21),
    .B2(_0424_),
    .C1(_0343_),
    .X(_0398_));
 sky130_fd_sc_hd__a211o_1 _1731_ (.A1(\phase_pwm_inst.counter[24] ),
    .A2(_0525_),
    .B1(_0397_),
    .C1(_0398_),
    .X(_0399_));
 sky130_fd_sc_hd__o31a_1 _1732_ (.A1(_0395_),
    .A2(_0396_),
    .A3(_0399_),
    .B1(_0348_),
    .X(_0400_));
 sky130_fd_sc_hd__o22a_1 _1733_ (.A1(_0421_),
    .A2(net25),
    .B1(_0339_),
    .B2(_0400_),
    .X(_0036_));
 sky130_fd_sc_hd__xor2_1 _1734_ (.A(\normal_mode_inst.timer_cnt[0] ),
    .B(\normal_mode_inst.timer_cnt[1] ),
    .X(_0049_));
 sky130_fd_sc_hd__a21oi_1 _1735_ (.A1(\normal_mode_inst.timer_cnt[0] ),
    .A2(\normal_mode_inst.timer_cnt[1] ),
    .B1(\normal_mode_inst.timer_cnt[2] ),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _1736_ (.A(_0762_),
    .B(_0401_),
    .Y(_0060_));
 sky130_fd_sc_hd__nor2_1 _1737_ (.A(\normal_mode_inst.timer_cnt[3] ),
    .B(_0762_),
    .Y(_0402_));
 sky130_fd_sc_hd__nor2_1 _1738_ (.A(_0763_),
    .B(_0402_),
    .Y(_0063_));
 sky130_fd_sc_hd__or2_1 _1739_ (.A(\normal_mode_inst.timer_cnt[4] ),
    .B(_0763_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _1740_ (.A(_0764_),
    .B(_0403_),
    .X(_0064_));
 sky130_fd_sc_hd__xnor2_1 _1741_ (.A(\normal_mode_inst.timer_cnt[5] ),
    .B(_0764_),
    .Y(_0065_));
 sky130_fd_sc_hd__a31o_1 _1742_ (.A1(\normal_mode_inst.timer_cnt[5] ),
    .A2(\normal_mode_inst.timer_cnt[4] ),
    .A3(_0763_),
    .B1(\normal_mode_inst.timer_cnt[6] ),
    .X(_0404_));
 sky130_fd_sc_hd__and2b_1 _1743_ (.A_N(_0765_),
    .B(_0404_),
    .X(_0066_));
 sky130_fd_sc_hd__or2_1 _1744_ (.A(\normal_mode_inst.timer_cnt[7] ),
    .B(_0765_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _1745_ (.A(_0766_),
    .B(_0405_),
    .X(_0067_));
 sky130_fd_sc_hd__xnor2_1 _1746_ (.A(\normal_mode_inst.timer_cnt[8] ),
    .B(_0766_),
    .Y(_0068_));
 sky130_fd_sc_hd__a31o_1 _1747_ (.A1(\normal_mode_inst.timer_cnt[7] ),
    .A2(\normal_mode_inst.timer_cnt[8] ),
    .A3(_0765_),
    .B1(\normal_mode_inst.timer_cnt[9] ),
    .X(_0406_));
 sky130_fd_sc_hd__and2b_1 _1748_ (.A_N(_0767_),
    .B(_0406_),
    .X(_0069_));
 sky130_fd_sc_hd__or2_1 _1749_ (.A(\normal_mode_inst.timer_cnt[10] ),
    .B(_0767_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _1750_ (.A(_0768_),
    .B(_0407_),
    .X(_0039_));
 sky130_fd_sc_hd__xnor2_1 _1751_ (.A(\normal_mode_inst.timer_cnt[11] ),
    .B(_0768_),
    .Y(_0040_));
 sky130_fd_sc_hd__a31o_1 _1752_ (.A1(\normal_mode_inst.timer_cnt[11] ),
    .A2(\normal_mode_inst.timer_cnt[10] ),
    .A3(_0767_),
    .B1(\normal_mode_inst.timer_cnt[12] ),
    .X(_0408_));
 sky130_fd_sc_hd__and2b_1 _1753_ (.A_N(_0769_),
    .B(_0408_),
    .X(_0041_));
 sky130_fd_sc_hd__or2_1 _1754_ (.A(\normal_mode_inst.timer_cnt[13] ),
    .B(_0769_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _1755_ (.A(_0770_),
    .B(_0409_),
    .X(_0042_));
 sky130_fd_sc_hd__xnor2_1 _1756_ (.A(\normal_mode_inst.timer_cnt[14] ),
    .B(_0770_),
    .Y(_0043_));
 sky130_fd_sc_hd__a31o_1 _1757_ (.A1(\normal_mode_inst.timer_cnt[13] ),
    .A2(\normal_mode_inst.timer_cnt[14] ),
    .A3(_0769_),
    .B1(\normal_mode_inst.timer_cnt[15] ),
    .X(_0410_));
 sky130_fd_sc_hd__and2b_1 _1758_ (.A_N(_0771_),
    .B(_0410_),
    .X(_0044_));
 sky130_fd_sc_hd__or2_1 _1759_ (.A(\normal_mode_inst.timer_cnt[16] ),
    .B(_0771_),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _1760_ (.A(_0772_),
    .B(_0411_),
    .X(_0045_));
 sky130_fd_sc_hd__xnor2_1 _1761_ (.A(\normal_mode_inst.timer_cnt[17] ),
    .B(_0772_),
    .Y(_0046_));
 sky130_fd_sc_hd__a31o_1 _1762_ (.A1(\normal_mode_inst.timer_cnt[17] ),
    .A2(\normal_mode_inst.timer_cnt[16] ),
    .A3(_0771_),
    .B1(\normal_mode_inst.timer_cnt[18] ),
    .X(_0412_));
 sky130_fd_sc_hd__and2b_1 _1763_ (.A_N(_0773_),
    .B(_0412_),
    .X(_0047_));
 sky130_fd_sc_hd__or2_1 _1764_ (.A(\normal_mode_inst.timer_cnt[19] ),
    .B(_0773_),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _1765_ (.A(_0774_),
    .B(_0413_),
    .X(_0048_));
 sky130_fd_sc_hd__xnor2_1 _1766_ (.A(\normal_mode_inst.timer_cnt[20] ),
    .B(_0774_),
    .Y(_0050_));
 sky130_fd_sc_hd__a31o_1 _1767_ (.A1(\normal_mode_inst.timer_cnt[19] ),
    .A2(\normal_mode_inst.timer_cnt[20] ),
    .A3(_0773_),
    .B1(\normal_mode_inst.timer_cnt[21] ),
    .X(_0414_));
 sky130_fd_sc_hd__and2b_1 _1768_ (.A_N(_0775_),
    .B(_0414_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _1769_ (.A(\normal_mode_inst.timer_cnt[22] ),
    .B(_0775_),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _1770_ (.A(_0776_),
    .B(_0415_),
    .X(_0052_));
 sky130_fd_sc_hd__xnor2_1 _1771_ (.A(\normal_mode_inst.timer_cnt[23] ),
    .B(_0776_),
    .Y(_0053_));
 sky130_fd_sc_hd__a31o_1 _1772_ (.A1(\normal_mode_inst.timer_cnt[23] ),
    .A2(\normal_mode_inst.timer_cnt[22] ),
    .A3(_0775_),
    .B1(\normal_mode_inst.timer_cnt[24] ),
    .X(_0416_));
 sky130_fd_sc_hd__and2b_1 _1773_ (.A_N(_0777_),
    .B(_0416_),
    .X(_0054_));
 sky130_fd_sc_hd__xor2_1 _1774_ (.A(\normal_mode_inst.timer_cnt[25] ),
    .B(_0777_),
    .X(_0055_));
 sky130_fd_sc_hd__a21oi_1 _1775_ (.A1(\normal_mode_inst.timer_cnt[25] ),
    .A2(_0777_),
    .B1(\normal_mode_inst.timer_cnt[26] ),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _1776_ (.A(_0778_),
    .B(_0417_),
    .Y(_0056_));
 sky130_fd_sc_hd__nor2_1 _1777_ (.A(\normal_mode_inst.timer_cnt[27] ),
    .B(_0778_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _1778_ (.A(_0779_),
    .B(_0418_),
    .Y(_0057_));
 sky130_fd_sc_hd__xor2_1 _1779_ (.A(\normal_mode_inst.timer_cnt[28] ),
    .B(_0779_),
    .X(_0058_));
 sky130_fd_sc_hd__a21oi_1 _1780_ (.A1(\normal_mode_inst.timer_cnt[28] ),
    .A2(_0779_),
    .B1(\normal_mode_inst.timer_cnt[29] ),
    .Y(_0419_));
 sky130_fd_sc_hd__nor2_1 _1781_ (.A(_0780_),
    .B(_0419_),
    .Y(_0059_));
 sky130_fd_sc_hd__xor2_1 _1782_ (.A(\normal_mode_inst.timer_cnt[30] ),
    .B(_0780_),
    .X(_0061_));
 sky130_fd_sc_hd__a21o_1 _1783_ (.A1(\normal_mode_inst.timer_cnt[30] ),
    .A2(_0780_),
    .B1(\normal_mode_inst.timer_cnt[31] ),
    .X(_0420_));
 sky130_fd_sc_hd__and2b_1 _1784_ (.A_N(_0034_),
    .B(_0420_),
    .X(_0062_));
 sky130_fd_sc_hd__nor3b_1 _1785_ (.A(net97),
    .B(net98),
    .C_N(irq_timer_normal),
    .Y(net102));
 sky130_fd_sc_hd__inv_2 _1786_ (.A(net99),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1787_ (.A(net99),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1788_ (.A(net99),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1789_ (.A(net99),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1790_ (.A(net99),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1791_ (.A(net99),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1792_ (.A(net99),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1793_ (.A(net99),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1794_ (.A(net99),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1795_ (.A(net99),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1796_ (.A(net99),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1797_ (.A(net99),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1798_ (.A(net99),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1799_ (.A(net99),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1800_ (.A(net99),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1801_ (.A(net99),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1802_ (.A(net99),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1803_ (.A(net99),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1804_ (.A(net99),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1805_ (.A(net99),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1806_ (.A(net99),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1807_ (.A(net99),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1808_ (.A(net99),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1809_ (.A(net99),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1810_ (.A(net99),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1811_ (.A(net99),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1812_ (.A(net99),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1813_ (.A(net99),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1814_ (.A(net99),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1815_ (.A(net99),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1816_ (.A(net99),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1817_ (.A(net99),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1818_ (.A(net99),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1819_ (.A(net99),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1820_ (.A(net99),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1821_ (.A(net99),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1822_ (.A(net99),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1823_ (.A(net99),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1824_ (.A(net99),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1825_ (.A(net99),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(net99),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(net99),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1828_ (.A(net99),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1829_ (.A(net99),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(net99),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1831_ (.A(net99),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1832_ (.A(net99),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(net99),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1834_ (.A(net99),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1835_ (.A(net99),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1836_ (.A(net99),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1837_ (.A(net99),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1838_ (.A(net99),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(net99),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(net99),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1841_ (.A(net99),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1842_ (.A(net99),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1843_ (.A(net99),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1844_ (.A(net99),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1845_ (.A(net99),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1846_ (.A(net99),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(net99),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1848_ (.A(net99),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1849_ (.A(net99),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(net99),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(net99),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(net99),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1853_ (.A(net99),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1854_ (.A(net99),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1855_ (.A(net99),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(net99),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1857_ (.A(net99),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1858_ (.A(net99),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(net99),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1860_ (.A(net99),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1861_ (.A(net99),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(net99),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1863_ (.A(net99),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1864_ (.A(net99),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1865_ (.A(net99),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1866_ (.A(net99),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1867_ (.A(net99),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(net99),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1869_ (.A(net99),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1870_ (.A(net99),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1871_ (.A(net99),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(net99),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(net99),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1874_ (.A(net99),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1875_ (.A(net99),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1876_ (.A(net99),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1877_ (.A(net99),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1878_ (.A(net99),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(net99),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1880_ (.A(net99),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1881_ (.A(net99),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1882_ (.A(net99),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1883_ (.A(net99),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1884_ (.A(net99),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1885_ (.A(net99),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1886_ (.A(net99),
    .Y(_0171_));
 sky130_fd_sc_hd__dfrtp_4 _1887_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0172_),
    .RESET_B(_0070_),
    .Q(\phase_pwm_inst.counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1888_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0173_),
    .RESET_B(_0071_),
    .Q(\phase_pwm_inst.counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1889_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0174_),
    .RESET_B(_0072_),
    .Q(\phase_pwm_inst.counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1890_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0175_),
    .RESET_B(_0073_),
    .Q(\phase_pwm_inst.counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1891_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0176_),
    .RESET_B(_0074_),
    .Q(\phase_pwm_inst.counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1892_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0177_),
    .RESET_B(_0075_),
    .Q(\phase_pwm_inst.counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1893_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0178_),
    .RESET_B(_0076_),
    .Q(\phase_pwm_inst.counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1894_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0179_),
    .RESET_B(_0077_),
    .Q(\phase_pwm_inst.counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _1895_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0180_),
    .RESET_B(_0078_),
    .Q(\phase_pwm_inst.counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1896_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0181_),
    .RESET_B(_0079_),
    .Q(\phase_pwm_inst.counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1897_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0182_),
    .RESET_B(_0080_),
    .Q(\phase_pwm_inst.counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _1898_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0183_),
    .RESET_B(_0081_),
    .Q(\phase_pwm_inst.counter[11] ));
 sky130_fd_sc_hd__dfrtp_4 _1899_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0184_),
    .RESET_B(_0082_),
    .Q(\phase_pwm_inst.counter[12] ));
 sky130_fd_sc_hd__dfrtp_4 _1900_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0185_),
    .RESET_B(_0083_),
    .Q(\phase_pwm_inst.counter[13] ));
 sky130_fd_sc_hd__dfrtp_4 _1901_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0186_),
    .RESET_B(_0084_),
    .Q(\phase_pwm_inst.counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _1902_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0187_),
    .RESET_B(_0085_),
    .Q(\phase_pwm_inst.counter[15] ));
 sky130_fd_sc_hd__dfrtp_4 _1903_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0188_),
    .RESET_B(_0086_),
    .Q(\phase_pwm_inst.counter[16] ));
 sky130_fd_sc_hd__dfrtp_4 _1904_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0189_),
    .RESET_B(_0087_),
    .Q(\phase_pwm_inst.counter[17] ));
 sky130_fd_sc_hd__dfrtp_4 _1905_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0190_),
    .RESET_B(_0088_),
    .Q(\phase_pwm_inst.counter[18] ));
 sky130_fd_sc_hd__dfrtp_4 _1906_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0191_),
    .RESET_B(_0089_),
    .Q(\phase_pwm_inst.counter[19] ));
 sky130_fd_sc_hd__dfrtp_4 _1907_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0192_),
    .RESET_B(_0090_),
    .Q(\phase_pwm_inst.counter[20] ));
 sky130_fd_sc_hd__dfrtp_2 _1908_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0193_),
    .RESET_B(_0091_),
    .Q(\phase_pwm_inst.counter[21] ));
 sky130_fd_sc_hd__dfrtp_4 _1909_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0194_),
    .RESET_B(_0092_),
    .Q(\phase_pwm_inst.counter[22] ));
 sky130_fd_sc_hd__dfrtp_4 _1910_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0195_),
    .RESET_B(_0093_),
    .Q(\phase_pwm_inst.counter[23] ));
 sky130_fd_sc_hd__dfrtp_4 _1911_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0196_),
    .RESET_B(_0094_),
    .Q(\phase_pwm_inst.counter[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1912_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0197_),
    .RESET_B(_0095_),
    .Q(\phase_pwm_inst.counter[25] ));
 sky130_fd_sc_hd__dfrtp_4 _1913_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0198_),
    .RESET_B(_0096_),
    .Q(\phase_pwm_inst.counter[26] ));
 sky130_fd_sc_hd__dfrtp_4 _1914_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0199_),
    .RESET_B(_0097_),
    .Q(\phase_pwm_inst.counter[27] ));
 sky130_fd_sc_hd__dfrtp_4 _1915_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0200_),
    .RESET_B(_0098_),
    .Q(\phase_pwm_inst.counter[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1916_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0201_),
    .RESET_B(_0099_),
    .Q(\phase_pwm_inst.counter[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1917_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0202_),
    .RESET_B(_0100_),
    .Q(\phase_pwm_inst.counter[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1918_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0203_),
    .RESET_B(_0101_),
    .Q(\phase_pwm_inst.counter[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1919_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0034_),
    .RESET_B(_0102_),
    .Q(irq_timer_normal));
 sky130_fd_sc_hd__dfrtp_1 _1920_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0038_),
    .RESET_B(_0103_),
    .Q(\normal_mode_inst.timer_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1921_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0049_),
    .RESET_B(_0104_),
    .Q(\normal_mode_inst.timer_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1922_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0060_),
    .RESET_B(_0105_),
    .Q(\normal_mode_inst.timer_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1923_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0063_),
    .RESET_B(_0106_),
    .Q(\normal_mode_inst.timer_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1924_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0064_),
    .RESET_B(_0107_),
    .Q(\normal_mode_inst.timer_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1925_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0065_),
    .RESET_B(_0108_),
    .Q(\normal_mode_inst.timer_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1926_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0066_),
    .RESET_B(_0109_),
    .Q(\normal_mode_inst.timer_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1927_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0067_),
    .RESET_B(_0110_),
    .Q(\normal_mode_inst.timer_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1928_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0068_),
    .RESET_B(_0111_),
    .Q(\normal_mode_inst.timer_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1929_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0069_),
    .RESET_B(_0112_),
    .Q(\normal_mode_inst.timer_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1930_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0039_),
    .RESET_B(_0113_),
    .Q(\normal_mode_inst.timer_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1931_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0040_),
    .RESET_B(_0114_),
    .Q(\normal_mode_inst.timer_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1932_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0041_),
    .RESET_B(_0115_),
    .Q(\normal_mode_inst.timer_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1933_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0042_),
    .RESET_B(_0116_),
    .Q(\normal_mode_inst.timer_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1934_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0043_),
    .RESET_B(_0117_),
    .Q(\normal_mode_inst.timer_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1935_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0044_),
    .RESET_B(_0118_),
    .Q(\normal_mode_inst.timer_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1936_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0045_),
    .RESET_B(_0119_),
    .Q(\normal_mode_inst.timer_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1937_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0046_),
    .RESET_B(_0120_),
    .Q(\normal_mode_inst.timer_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1938_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0047_),
    .RESET_B(_0121_),
    .Q(\normal_mode_inst.timer_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_1 _1939_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0048_),
    .RESET_B(_0122_),
    .Q(\normal_mode_inst.timer_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_1 _1940_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0050_),
    .RESET_B(_0123_),
    .Q(\normal_mode_inst.timer_cnt[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1941_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0051_),
    .RESET_B(_0124_),
    .Q(\normal_mode_inst.timer_cnt[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1942_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0052_),
    .RESET_B(_0125_),
    .Q(\normal_mode_inst.timer_cnt[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1943_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0053_),
    .RESET_B(_0126_),
    .Q(\normal_mode_inst.timer_cnt[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1944_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0054_),
    .RESET_B(_0127_),
    .Q(\normal_mode_inst.timer_cnt[24] ));
 sky130_fd_sc_hd__dfrtp_1 _1945_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0055_),
    .RESET_B(_0128_),
    .Q(\normal_mode_inst.timer_cnt[25] ));
 sky130_fd_sc_hd__dfrtp_1 _1946_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0056_),
    .RESET_B(_0129_),
    .Q(\normal_mode_inst.timer_cnt[26] ));
 sky130_fd_sc_hd__dfrtp_1 _1947_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0057_),
    .RESET_B(_0130_),
    .Q(\normal_mode_inst.timer_cnt[27] ));
 sky130_fd_sc_hd__dfrtp_1 _1948_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0058_),
    .RESET_B(_0131_),
    .Q(\normal_mode_inst.timer_cnt[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1949_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0059_),
    .RESET_B(_0132_),
    .Q(\normal_mode_inst.timer_cnt[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1950_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0061_),
    .RESET_B(_0133_),
    .Q(\normal_mode_inst.timer_cnt[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1951_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0062_),
    .RESET_B(_0134_),
    .Q(\normal_mode_inst.timer_cnt[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1952_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0033_),
    .RESET_B(_0135_),
    .Q(\fast_pwm_inst.pwm_outb ));
 sky130_fd_sc_hd__dfrtp_1 _1953_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0032_),
    .RESET_B(_0136_),
    .Q(\fast_pwm_inst.pwm_outa ));
 sky130_fd_sc_hd__dfrtp_1 _1954_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0000_),
    .RESET_B(_0137_),
    .Q(\fast_pwm_inst.pwm_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1955_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0011_),
    .RESET_B(_0138_),
    .Q(\fast_pwm_inst.pwm_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1956_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0022_),
    .RESET_B(_0139_),
    .Q(\fast_pwm_inst.pwm_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1957_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0025_),
    .RESET_B(_0140_),
    .Q(\fast_pwm_inst.pwm_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1958_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0026_),
    .RESET_B(_0141_),
    .Q(\fast_pwm_inst.pwm_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1959_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0027_),
    .RESET_B(_0142_),
    .Q(\fast_pwm_inst.pwm_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1960_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0028_),
    .RESET_B(_0143_),
    .Q(\fast_pwm_inst.pwm_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1961_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0029_),
    .RESET_B(_0144_),
    .Q(\fast_pwm_inst.pwm_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1962_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0030_),
    .RESET_B(_0145_),
    .Q(\fast_pwm_inst.pwm_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1963_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0031_),
    .RESET_B(_0146_),
    .Q(\fast_pwm_inst.pwm_counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _1964_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0001_),
    .RESET_B(_0147_),
    .Q(\fast_pwm_inst.pwm_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1965_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0002_),
    .RESET_B(_0148_),
    .Q(\fast_pwm_inst.pwm_counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 _1966_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0003_),
    .RESET_B(_0149_),
    .Q(\fast_pwm_inst.pwm_counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 _1967_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0004_),
    .RESET_B(_0150_),
    .Q(\fast_pwm_inst.pwm_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1968_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0005_),
    .RESET_B(_0151_),
    .Q(\fast_pwm_inst.pwm_counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _1969_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0006_),
    .RESET_B(_0152_),
    .Q(\fast_pwm_inst.pwm_counter[15] ));
 sky130_fd_sc_hd__dfrtp_2 _1970_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0007_),
    .RESET_B(_0153_),
    .Q(\fast_pwm_inst.pwm_counter[16] ));
 sky130_fd_sc_hd__dfrtp_1 _1971_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0008_),
    .RESET_B(_0154_),
    .Q(\fast_pwm_inst.pwm_counter[17] ));
 sky130_fd_sc_hd__dfrtp_1 _1972_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0009_),
    .RESET_B(_0155_),
    .Q(\fast_pwm_inst.pwm_counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 _1973_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0010_),
    .RESET_B(_0156_),
    .Q(\fast_pwm_inst.pwm_counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 _1974_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0012_),
    .RESET_B(_0157_),
    .Q(\fast_pwm_inst.pwm_counter[20] ));
 sky130_fd_sc_hd__dfrtp_4 _1975_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0013_),
    .RESET_B(_0158_),
    .Q(\fast_pwm_inst.pwm_counter[21] ));
 sky130_fd_sc_hd__dfrtp_4 _1976_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0014_),
    .RESET_B(_0159_),
    .Q(\fast_pwm_inst.pwm_counter[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1977_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0015_),
    .RESET_B(_0160_),
    .Q(\fast_pwm_inst.pwm_counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 _1978_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0016_),
    .RESET_B(_0161_),
    .Q(\fast_pwm_inst.pwm_counter[24] ));
 sky130_fd_sc_hd__dfrtp_4 _1979_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0017_),
    .RESET_B(_0162_),
    .Q(\fast_pwm_inst.pwm_counter[25] ));
 sky130_fd_sc_hd__dfrtp_2 _1980_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0018_),
    .RESET_B(_0163_),
    .Q(\fast_pwm_inst.pwm_counter[26] ));
 sky130_fd_sc_hd__dfrtp_2 _1981_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0019_),
    .RESET_B(_0164_),
    .Q(\fast_pwm_inst.pwm_counter[27] ));
 sky130_fd_sc_hd__dfrtp_4 _1982_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0020_),
    .RESET_B(_0165_),
    .Q(\fast_pwm_inst.pwm_counter[28] ));
 sky130_fd_sc_hd__dfrtp_2 _1983_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0021_),
    .RESET_B(_0166_),
    .Q(\fast_pwm_inst.pwm_counter[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1984_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0023_),
    .RESET_B(_0167_),
    .Q(\fast_pwm_inst.pwm_counter[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1985_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0024_),
    .RESET_B(_0168_),
    .Q(\fast_pwm_inst.pwm_counter[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1986_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0037_),
    .RESET_B(_0169_),
    .Q(\phase_pwm_inst.pwm_outb ));
 sky130_fd_sc_hd__dfrtp_1 _1987_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0036_),
    .RESET_B(_0170_),
    .Q(\phase_pwm_inst.pwm_outa ));
 sky130_fd_sc_hd__dfrtp_4 _1988_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0035_),
    .RESET_B(_0171_),
    .Q(\phase_pwm_inst.direction ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_373 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(PWM_CNTA[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(PWM_CNTA[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(PWM_CNTA[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(PWM_CNTA[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(PWM_CNTA[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(PWM_CNTA[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(PWM_CNTA[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(PWM_CNTA[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(PWM_CNTA[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(PWM_CNTA[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(PWM_CNTA[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(PWM_CNTA[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(PWM_CNTA[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(PWM_CNTA[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(PWM_CNTA[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(PWM_CNTA[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(PWM_CNTA[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(PWM_CNTA[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(PWM_CNTA[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(PWM_CNTA[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(PWM_CNTA[28]),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input22 (.A(PWM_CNTA[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(PWM_CNTA[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(PWM_CNTA[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(PWM_CNTA[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(PWM_CNTA[3]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(PWM_CNTA[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(PWM_CNTA[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(PWM_CNTA[6]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(PWM_CNTA[7]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(PWM_CNTA[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(PWM_CNTA[9]),
    .X(net32));
 sky130_fd_sc_hd__dlymetal6s2s_1 input33 (.A(PWM_CNTB[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(PWM_CNTB[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(PWM_CNTB[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(PWM_CNTB[12]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(PWM_CNTB[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(PWM_CNTB[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(PWM_CNTB[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(PWM_CNTB[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(PWM_CNTB[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(PWM_CNTB[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(PWM_CNTB[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(PWM_CNTB[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(PWM_CNTB[20]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input46 (.A(PWM_CNTB[21]),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 input47 (.A(PWM_CNTB[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(PWM_CNTB[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(PWM_CNTB[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(PWM_CNTB[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(PWM_CNTB[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(PWM_CNTB[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(PWM_CNTB[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(PWM_CNTB[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(PWM_CNTB[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(PWM_CNTB[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(PWM_CNTB[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 input58 (.A(PWM_CNTB[3]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(PWM_CNTB[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(PWM_CNTB[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(PWM_CNTB[6]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(PWM_CNTB[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(PWM_CNTB[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input64 (.A(PWM_CNTB[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(TIMER_TOP[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(TIMER_TOP[10]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(TIMER_TOP[11]),
    .X(net67));
 sky130_fd_sc_hd__dlymetal6s2s_1 input68 (.A(TIMER_TOP[12]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(TIMER_TOP[13]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(TIMER_TOP[14]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(TIMER_TOP[15]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(TIMER_TOP[16]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(TIMER_TOP[17]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(TIMER_TOP[18]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(TIMER_TOP[19]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(TIMER_TOP[1]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 input77 (.A(TIMER_TOP[20]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(TIMER_TOP[21]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(TIMER_TOP[22]),
    .X(net79));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(TIMER_TOP[23]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(TIMER_TOP[24]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(TIMER_TOP[25]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(TIMER_TOP[26]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(TIMER_TOP[27]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(TIMER_TOP[28]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(TIMER_TOP[29]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(TIMER_TOP[2]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_2 input88 (.A(TIMER_TOP[30]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(TIMER_TOP[31]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(TIMER_TOP[3]),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input91 (.A(TIMER_TOP[4]),
    .X(net91));
 sky130_fd_sc_hd__dlymetal6s2s_1 input92 (.A(TIMER_TOP[5]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(TIMER_TOP[6]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 input94 (.A(TIMER_TOP[7]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(TIMER_TOP[8]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input96 (.A(TIMER_TOP[9]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(TMR_MODE[0]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(TMR_MODE[1]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_16 input99 (.A(reset),
    .X(net99));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(PWM_OUTA));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(PWM_OUTB));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(timer_interrupt));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload6 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net100));
 sky130_fd_sc_hd__decap_8 FILLER_0_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
endmodule
