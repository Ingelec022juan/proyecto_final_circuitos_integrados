VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Timer_PWM_Generator
  CLASS BLOCK ;
  FOREIGN Timer_PWM_Generator ;
  ORIGIN 0.000 0.000 ;
  SIZE 154.515 BY 165.235 ;
  PIN PWM_CNTA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 161.235 42.230 165.235 ;
    END
  END PWM_CNTA[0]
  PIN PWM_CNTA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END PWM_CNTA[10]
  PIN PWM_CNTA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END PWM_CNTA[11]
  PIN PWM_CNTA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 161.235 77.650 165.235 ;
    END
  END PWM_CNTA[12]
  PIN PWM_CNTA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END PWM_CNTA[13]
  PIN PWM_CNTA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 61.240 154.515 61.840 ;
    END
  END PWM_CNTA[14]
  PIN PWM_CNTA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END PWM_CNTA[15]
  PIN PWM_CNTA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 96.690 161.235 96.970 165.235 ;
    END
  END PWM_CNTA[16]
  PIN PWM_CNTA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END PWM_CNTA[17]
  PIN PWM_CNTA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END PWM_CNTA[18]
  PIN PWM_CNTA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 129.240 154.515 129.840 ;
    END
  END PWM_CNTA[19]
  PIN PWM_CNTA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END PWM_CNTA[1]
  PIN PWM_CNTA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END PWM_CNTA[20]
  PIN PWM_CNTA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 37.440 154.515 38.040 ;
    END
  END PWM_CNTA[21]
  PIN PWM_CNTA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END PWM_CNTA[22]
  PIN PWM_CNTA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 85.040 154.515 85.640 ;
    END
  END PWM_CNTA[23]
  PIN PWM_CNTA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END PWM_CNTA[24]
  PIN PWM_CNTA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END PWM_CNTA[25]
  PIN PWM_CNTA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 132.110 161.235 132.390 165.235 ;
    END
  END PWM_CNTA[26]
  PIN PWM_CNTA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END PWM_CNTA[27]
  PIN PWM_CNTA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 30.640 154.515 31.240 ;
    END
  END PWM_CNTA[28]
  PIN PWM_CNTA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 91.840 154.515 92.440 ;
    END
  END PWM_CNTA[29]
  PIN PWM_CNTA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 149.640 154.515 150.240 ;
    END
  END PWM_CNTA[2]
  PIN PWM_CNTA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 161.235 13.250 165.235 ;
    END
  END PWM_CNTA[30]
  PIN PWM_CNTA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END PWM_CNTA[31]
  PIN PWM_CNTA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.570 161.235 109.850 165.235 ;
    END
  END PWM_CNTA[3]
  PIN PWM_CNTA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END PWM_CNTA[4]
  PIN PWM_CNTA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 161.235 145.270 165.235 ;
    END
  END PWM_CNTA[5]
  PIN PWM_CNTA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 156.440 154.515 157.040 ;
    END
  END PWM_CNTA[6]
  PIN PWM_CNTA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END PWM_CNTA[7]
  PIN PWM_CNTA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END PWM_CNTA[8]
  PIN PWM_CNTA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END PWM_CNTA[9]
  PIN PWM_CNTB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 163.240 154.515 163.840 ;
    END
  END PWM_CNTB[0]
  PIN PWM_CNTB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 125.670 161.235 125.950 165.235 ;
    END
  END PWM_CNTB[10]
  PIN PWM_CNTB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 10.240 154.515 10.840 ;
    END
  END PWM_CNTB[11]
  PIN PWM_CNTB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END PWM_CNTB[12]
  PIN PWM_CNTB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 74.840 154.515 75.440 ;
    END
  END PWM_CNTB[13]
  PIN PWM_CNTB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 54.440 154.515 55.040 ;
    END
  END PWM_CNTB[14]
  PIN PWM_CNTB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 161.235 48.670 165.235 ;
    END
  END PWM_CNTB[15]
  PIN PWM_CNTB[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 161.235 55.110 165.235 ;
    END
  END PWM_CNTB[16]
  PIN PWM_CNTB[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 122.440 154.515 123.040 ;
    END
  END PWM_CNTB[17]
  PIN PWM_CNTB[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END PWM_CNTB[18]
  PIN PWM_CNTB[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END PWM_CNTB[19]
  PIN PWM_CNTB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 136.040 154.515 136.640 ;
    END
  END PWM_CNTB[1]
  PIN PWM_CNTB[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 3.440 154.515 4.040 ;
    END
  END PWM_CNTB[20]
  PIN PWM_CNTB[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 161.235 84.090 165.235 ;
    END
  END PWM_CNTB[21]
  PIN PWM_CNTB[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END PWM_CNTB[22]
  PIN PWM_CNTB[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 161.235 35.790 165.235 ;
    END
  END PWM_CNTB[23]
  PIN PWM_CNTB[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 161.235 61.550 165.235 ;
    END
  END PWM_CNTB[24]
  PIN PWM_CNTB[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 142.840 154.515 143.440 ;
    END
  END PWM_CNTB[25]
  PIN PWM_CNTB[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 0.040 154.515 0.640 ;
    END
  END PWM_CNTB[26]
  PIN PWM_CNTB[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 161.235 74.430 165.235 ;
    END
  END PWM_CNTB[27]
  PIN PWM_CNTB[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END PWM_CNTB[28]
  PIN PWM_CNTB[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 40.840 154.515 41.440 ;
    END
  END PWM_CNTB[29]
  PIN PWM_CNTB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 105.440 154.515 106.040 ;
    END
  END PWM_CNTB[2]
  PIN PWM_CNTB[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END PWM_CNTB[30]
  PIN PWM_CNTB[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 161.235 90.530 165.235 ;
    END
  END PWM_CNTB[31]
  PIN PWM_CNTB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 161.235 26.130 165.235 ;
    END
  END PWM_CNTB[3]
  PIN PWM_CNTB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END PWM_CNTB[4]
  PIN PWM_CNTB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END PWM_CNTB[5]
  PIN PWM_CNTB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END PWM_CNTB[6]
  PIN PWM_CNTB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END PWM_CNTB[7]
  PIN PWM_CNTB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END PWM_CNTB[8]
  PIN PWM_CNTB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END PWM_CNTB[9]
  PIN PWM_OUTA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END PWM_OUTA
  PIN PWM_OUTB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 150.515 47.640 154.515 48.240 ;
    END
  END PWM_OUTB
  PIN TIMER_TOP[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END TIMER_TOP[0]
  PIN TIMER_TOP[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END TIMER_TOP[10]
  PIN TIMER_TOP[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 17.040 154.515 17.640 ;
    END
  END TIMER_TOP[11]
  PIN TIMER_TOP[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END TIMER_TOP[12]
  PIN TIMER_TOP[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 68.040 154.515 68.640 ;
    END
  END TIMER_TOP[13]
  PIN TIMER_TOP[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 112.240 154.515 112.840 ;
    END
  END TIMER_TOP[14]
  PIN TIMER_TOP[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END TIMER_TOP[15]
  PIN TIMER_TOP[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 119.040 154.515 119.640 ;
    END
  END TIMER_TOP[16]
  PIN TIMER_TOP[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END TIMER_TOP[17]
  PIN TIMER_TOP[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END TIMER_TOP[18]
  PIN TIMER_TOP[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END TIMER_TOP[19]
  PIN TIMER_TOP[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END TIMER_TOP[1]
  PIN TIMER_TOP[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END TIMER_TOP[20]
  PIN TIMER_TOP[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 161.235 19.690 165.235 ;
    END
  END TIMER_TOP[21]
  PIN TIMER_TOP[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 161.235 67.990 165.235 ;
    END
  END TIMER_TOP[22]
  PIN TIMER_TOP[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END TIMER_TOP[23]
  PIN TIMER_TOP[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END TIMER_TOP[24]
  PIN TIMER_TOP[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END TIMER_TOP[25]
  PIN TIMER_TOP[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END TIMER_TOP[26]
  PIN TIMER_TOP[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.550 161.235 138.830 165.235 ;
    END
  END TIMER_TOP[27]
  PIN TIMER_TOP[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.130 161.235 103.410 165.235 ;
    END
  END TIMER_TOP[28]
  PIN TIMER_TOP[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END TIMER_TOP[29]
  PIN TIMER_TOP[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 161.235 151.710 165.235 ;
    END
  END TIMER_TOP[2]
  PIN TIMER_TOP[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 23.840 154.515 24.440 ;
    END
  END TIMER_TOP[30]
  PIN TIMER_TOP[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 161.235 0.370 165.235 ;
    END
  END TIMER_TOP[31]
  PIN TIMER_TOP[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END TIMER_TOP[3]
  PIN TIMER_TOP[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END TIMER_TOP[4]
  PIN TIMER_TOP[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END TIMER_TOP[5]
  PIN TIMER_TOP[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END TIMER_TOP[6]
  PIN TIMER_TOP[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 150.515 98.640 154.515 99.240 ;
    END
  END TIMER_TOP[7]
  PIN TIMER_TOP[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END TIMER_TOP[8]
  PIN TIMER_TOP[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 119.230 161.235 119.510 165.235 ;
    END
  END TIMER_TOP[9]
  PIN TMR_MODE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 161.235 113.070 165.235 ;
    END
  END TMR_MODE[0]
  PIN TMR_MODE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 6.530 161.235 6.810 165.235 ;
    END
  END TMR_MODE[1]
  PIN TMR_SRC[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 161.235 32.570 165.235 ;
    END
  END TMR_SRC[0]
  PIN TMR_SRC[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END TMR_SRC[1]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 152.560 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 152.560 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END reset
  PIN timer_interrupt
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 150.515 81.640 154.515 82.240 ;
    END
  END timer_interrupt
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 148.770 152.405 ;
      LAYER li1 ;
        RECT 5.520 10.795 148.580 152.405 ;
      LAYER met1 ;
        RECT 0.070 8.200 151.730 152.560 ;
      LAYER met2 ;
        RECT 0.650 160.955 6.250 163.725 ;
        RECT 7.090 160.955 12.690 163.725 ;
        RECT 13.530 160.955 19.130 163.725 ;
        RECT 19.970 160.955 25.570 163.725 ;
        RECT 26.410 160.955 32.010 163.725 ;
        RECT 32.850 160.955 35.230 163.725 ;
        RECT 36.070 160.955 41.670 163.725 ;
        RECT 42.510 160.955 48.110 163.725 ;
        RECT 48.950 160.955 54.550 163.725 ;
        RECT 55.390 160.955 60.990 163.725 ;
        RECT 61.830 160.955 67.430 163.725 ;
        RECT 68.270 160.955 73.870 163.725 ;
        RECT 74.710 160.955 77.090 163.725 ;
        RECT 77.930 160.955 83.530 163.725 ;
        RECT 84.370 160.955 89.970 163.725 ;
        RECT 90.810 160.955 96.410 163.725 ;
        RECT 97.250 160.955 102.850 163.725 ;
        RECT 103.690 160.955 109.290 163.725 ;
        RECT 110.130 160.955 112.510 163.725 ;
        RECT 113.350 160.955 118.950 163.725 ;
        RECT 119.790 160.955 125.390 163.725 ;
        RECT 126.230 160.955 131.830 163.725 ;
        RECT 132.670 160.955 138.270 163.725 ;
        RECT 139.110 160.955 144.710 163.725 ;
        RECT 145.550 160.955 151.150 163.725 ;
        RECT 0.100 4.280 151.700 160.955 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 9.470 4.280 ;
        RECT 10.310 0.155 15.910 4.280 ;
        RECT 16.750 0.155 22.350 4.280 ;
        RECT 23.190 0.155 28.790 4.280 ;
        RECT 29.630 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 51.330 4.280 ;
        RECT 52.170 0.155 57.770 4.280 ;
        RECT 58.610 0.155 64.210 4.280 ;
        RECT 65.050 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 86.750 4.280 ;
        RECT 87.590 0.155 93.190 4.280 ;
        RECT 94.030 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 128.610 4.280 ;
        RECT 129.450 0.155 135.050 4.280 ;
        RECT 135.890 0.155 141.490 4.280 ;
        RECT 142.330 0.155 147.930 4.280 ;
        RECT 148.770 0.155 151.700 4.280 ;
      LAYER met3 ;
        RECT 4.400 162.840 150.115 163.705 ;
        RECT 3.990 157.440 150.515 162.840 ;
        RECT 4.400 156.040 150.115 157.440 ;
        RECT 3.990 150.640 150.515 156.040 ;
        RECT 4.400 149.240 150.115 150.640 ;
        RECT 3.990 143.840 150.515 149.240 ;
        RECT 4.400 142.440 150.115 143.840 ;
        RECT 3.990 137.040 150.515 142.440 ;
        RECT 4.400 135.640 150.115 137.040 ;
        RECT 3.990 130.240 150.515 135.640 ;
        RECT 4.400 128.840 150.115 130.240 ;
        RECT 3.990 123.440 150.515 128.840 ;
        RECT 4.400 122.040 150.115 123.440 ;
        RECT 3.990 120.040 150.515 122.040 ;
        RECT 4.400 118.640 150.115 120.040 ;
        RECT 3.990 113.240 150.515 118.640 ;
        RECT 4.400 111.840 150.115 113.240 ;
        RECT 3.990 106.440 150.515 111.840 ;
        RECT 4.400 105.040 150.115 106.440 ;
        RECT 3.990 99.640 150.515 105.040 ;
        RECT 4.400 98.240 150.115 99.640 ;
        RECT 3.990 92.840 150.515 98.240 ;
        RECT 4.400 91.440 150.115 92.840 ;
        RECT 3.990 86.040 150.515 91.440 ;
        RECT 4.400 84.640 150.115 86.040 ;
        RECT 3.990 82.640 150.515 84.640 ;
        RECT 4.400 81.240 150.115 82.640 ;
        RECT 3.990 75.840 150.515 81.240 ;
        RECT 4.400 74.440 150.115 75.840 ;
        RECT 3.990 69.040 150.515 74.440 ;
        RECT 4.400 67.640 150.115 69.040 ;
        RECT 3.990 62.240 150.515 67.640 ;
        RECT 4.400 60.840 150.115 62.240 ;
        RECT 3.990 55.440 150.515 60.840 ;
        RECT 4.400 54.040 150.115 55.440 ;
        RECT 3.990 48.640 150.515 54.040 ;
        RECT 4.400 47.240 150.115 48.640 ;
        RECT 3.990 41.840 150.515 47.240 ;
        RECT 4.400 40.440 150.115 41.840 ;
        RECT 3.990 38.440 150.515 40.440 ;
        RECT 4.400 37.040 150.115 38.440 ;
        RECT 3.990 31.640 150.515 37.040 ;
        RECT 4.400 30.240 150.115 31.640 ;
        RECT 3.990 24.840 150.515 30.240 ;
        RECT 4.400 23.440 150.115 24.840 ;
        RECT 3.990 18.040 150.515 23.440 ;
        RECT 4.400 16.640 150.115 18.040 ;
        RECT 3.990 11.240 150.515 16.640 ;
        RECT 4.400 9.840 150.115 11.240 ;
        RECT 3.990 4.440 150.515 9.840 ;
        RECT 4.400 3.040 150.115 4.440 ;
        RECT 3.990 1.040 150.515 3.040 ;
        RECT 3.990 0.175 150.115 1.040 ;
      LAYER met4 ;
        RECT 30.655 11.055 88.945 145.345 ;
  END
END Timer_PWM_Generator
END LIBRARY

