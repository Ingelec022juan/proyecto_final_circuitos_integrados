magic
tech sky130A
magscale 1 2
timestamp 1732234192
<< viali >>
rect 2421 30277 2455 30311
rect 2789 30277 2823 30311
rect 8585 30277 8619 30311
rect 9873 30277 9907 30311
rect 15761 30277 15795 30311
rect 19625 30277 19659 30311
rect 20913 30277 20947 30311
rect 22109 30277 22143 30311
rect 25421 30277 25455 30311
rect 28089 30277 28123 30311
rect 3157 30209 3191 30243
rect 3985 30209 4019 30243
rect 5273 30209 5307 30243
rect 7205 30209 7239 30243
rect 11069 30209 11103 30243
rect 12357 30209 12391 30243
rect 13829 30209 13863 30243
rect 14933 30209 14967 30243
rect 16865 30209 16899 30243
rect 18153 30209 18187 30243
rect 22661 30209 22695 30243
rect 23949 30209 23983 30243
rect 26985 30209 27019 30243
rect 28457 30209 28491 30243
rect 29377 30209 29411 30243
rect 1409 30141 1443 30175
rect 1685 30141 1719 30175
rect 17141 30141 17175 30175
rect 27261 30141 27295 30175
rect 29101 30141 29135 30175
rect 2605 30073 2639 30107
rect 2973 30073 3007 30107
rect 3341 30073 3375 30107
rect 7389 30073 7423 30107
rect 8769 30073 8803 30107
rect 10057 30073 10091 30107
rect 20729 30073 20763 30107
rect 22293 30073 22327 30107
rect 27905 30073 27939 30107
rect 4169 30005 4203 30039
rect 5457 30005 5491 30039
rect 11253 30005 11287 30039
rect 12541 30005 12575 30039
rect 13645 30005 13679 30039
rect 15117 30005 15151 30039
rect 15669 30005 15703 30039
rect 18337 30005 18371 30039
rect 19533 30005 19567 30039
rect 22845 30005 22879 30039
rect 24133 30005 24167 30039
rect 25329 30005 25363 30039
rect 28273 30005 28307 30039
rect 1409 29665 1443 29699
rect 1685 29597 1719 29631
rect 13553 29597 13587 29631
rect 28549 29597 28583 29631
rect 28917 29597 28951 29631
rect 29285 29597 29319 29631
rect 2421 29529 2455 29563
rect 2605 29529 2639 29563
rect 28365 29529 28399 29563
rect 28733 29529 28767 29563
rect 13461 29461 13495 29495
rect 29193 29461 29227 29495
rect 19533 29257 19567 29291
rect 1409 29121 1443 29155
rect 11161 29121 11195 29155
rect 23121 29121 23155 29155
rect 29285 29121 29319 29155
rect 3157 29053 3191 29087
rect 14473 29053 14507 29087
rect 16497 29053 16531 29087
rect 17785 29053 17819 29087
rect 18061 29053 18095 29087
rect 11253 28985 11287 29019
rect 23213 28985 23247 29019
rect 29101 28985 29135 29019
rect 14730 28917 14764 28951
rect 15669 28713 15703 28747
rect 18889 28713 18923 28747
rect 8125 28645 8159 28679
rect 25789 28645 25823 28679
rect 12173 28577 12207 28611
rect 17233 28577 17267 28611
rect 19993 28577 20027 28611
rect 22201 28577 22235 28611
rect 22477 28577 22511 28611
rect 24133 28577 24167 28611
rect 7297 28509 7331 28543
rect 7481 28509 7515 28543
rect 7573 28509 7607 28543
rect 7665 28509 7699 28543
rect 8217 28509 8251 28543
rect 9137 28509 9171 28543
rect 10149 28509 10183 28543
rect 12449 28509 12483 28543
rect 12633 28509 12667 28543
rect 12725 28509 12759 28543
rect 12817 28509 12851 28543
rect 13645 28509 13679 28543
rect 15761 28509 15795 28543
rect 17417 28509 17451 28543
rect 17693 28509 17727 28543
rect 17885 28509 17919 28543
rect 18797 28509 18831 28543
rect 24041 28509 24075 28543
rect 24225 28509 24259 28543
rect 25513 28509 25547 28543
rect 27077 28509 27111 28543
rect 29101 28509 29135 28543
rect 10425 28441 10459 28475
rect 20269 28441 20303 28475
rect 22017 28441 22051 28475
rect 25789 28441 25823 28475
rect 27353 28441 27387 28475
rect 29009 28441 29043 28475
rect 7941 28373 7975 28407
rect 9045 28373 9079 28407
rect 13093 28373 13127 28407
rect 13737 28373 13771 28407
rect 17601 28373 17635 28407
rect 18061 28373 18095 28407
rect 23949 28373 23983 28407
rect 25605 28373 25639 28407
rect 28825 28373 28859 28407
rect 10517 28169 10551 28203
rect 11069 28169 11103 28203
rect 14381 28169 14415 28203
rect 14565 28169 14599 28203
rect 15501 28169 15535 28203
rect 15669 28169 15703 28203
rect 19073 28169 19107 28203
rect 19825 28169 19859 28203
rect 19993 28169 20027 28203
rect 21189 28169 21223 28203
rect 24501 28169 24535 28203
rect 8033 28101 8067 28135
rect 12909 28101 12943 28135
rect 14749 28101 14783 28135
rect 15301 28101 15335 28135
rect 16129 28101 16163 28135
rect 19165 28101 19199 28135
rect 19625 28101 19659 28135
rect 26709 28101 26743 28135
rect 5825 28033 5859 28067
rect 6377 28033 6411 28067
rect 6561 28033 6595 28067
rect 9873 28033 9907 28067
rect 10057 28033 10091 28067
rect 10149 28033 10183 28067
rect 10241 28033 10275 28067
rect 10701 28033 10735 28067
rect 10885 28033 10919 28067
rect 10977 28033 11011 28067
rect 11161 28033 11195 28067
rect 12633 28033 12667 28067
rect 15761 28033 15795 28067
rect 18521 28033 18555 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 19349 28033 19383 28067
rect 21281 28033 21315 28067
rect 23489 28033 23523 28067
rect 24133 28033 24167 28067
rect 24225 28033 24259 28067
rect 24409 28033 24443 28067
rect 24593 28033 24627 28067
rect 26801 28033 26835 28067
rect 27169 28033 27203 28067
rect 7757 27965 7791 27999
rect 9781 27965 9815 27999
rect 18245 27965 18279 27999
rect 23581 27965 23615 27999
rect 23949 27965 23983 27999
rect 24777 27965 24811 27999
rect 25053 27965 25087 27999
rect 26525 27965 26559 27999
rect 27077 27965 27111 27999
rect 27537 27965 27571 27999
rect 15117 27897 15151 27931
rect 16313 27897 16347 27931
rect 5917 27829 5951 27863
rect 6469 27829 6503 27863
rect 10793 27829 10827 27863
rect 14749 27829 14783 27863
rect 15485 27829 15519 27863
rect 16129 27829 16163 27863
rect 16773 27829 16807 27863
rect 19533 27829 19567 27863
rect 19809 27829 19843 27863
rect 23857 27829 23891 27863
rect 7297 27625 7331 27659
rect 8309 27625 8343 27659
rect 9965 27625 9999 27659
rect 11069 27625 11103 27659
rect 14197 27625 14231 27659
rect 14841 27625 14875 27659
rect 15853 27625 15887 27659
rect 17877 27625 17911 27659
rect 18061 27625 18095 27659
rect 18889 27625 18923 27659
rect 19901 27625 19935 27659
rect 23599 27625 23633 27659
rect 25329 27625 25363 27659
rect 25789 27625 25823 27659
rect 6561 27557 6595 27591
rect 10701 27557 10735 27591
rect 13185 27557 13219 27591
rect 17049 27557 17083 27591
rect 17509 27557 17543 27591
rect 19073 27557 19107 27591
rect 19533 27557 19567 27591
rect 4813 27489 4847 27523
rect 8033 27489 8067 27523
rect 20177 27489 20211 27523
rect 22109 27489 22143 27523
rect 1409 27421 1443 27455
rect 1685 27421 1719 27455
rect 7205 27421 7239 27455
rect 7389 27421 7423 27455
rect 7481 27421 7515 27455
rect 7757 27421 7791 27455
rect 8677 27421 8711 27455
rect 9137 27421 9171 27455
rect 9873 27421 9907 27455
rect 10057 27421 10091 27455
rect 11345 27421 11379 27455
rect 13553 27421 13587 27455
rect 14197 27421 14231 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 15117 27421 15151 27455
rect 15485 27421 15519 27455
rect 16957 27421 16991 27455
rect 19257 27421 19291 27455
rect 19441 27421 19475 27455
rect 23857 27421 23891 27455
rect 25145 27421 25179 27455
rect 25329 27421 25363 27455
rect 27629 27421 27663 27455
rect 5089 27353 5123 27387
rect 6929 27353 6963 27387
rect 7113 27353 7147 27387
rect 7849 27353 7883 27387
rect 8309 27353 8343 27387
rect 11069 27353 11103 27387
rect 11621 27353 11655 27387
rect 13737 27353 13771 27387
rect 14657 27353 14691 27387
rect 15669 27353 15703 27387
rect 17877 27353 17911 27387
rect 18705 27353 18739 27387
rect 18905 27353 18939 27387
rect 20453 27353 20487 27387
rect 25757 27353 25791 27387
rect 25973 27353 26007 27387
rect 27905 27353 27939 27387
rect 6745 27285 6779 27319
rect 7665 27285 7699 27319
rect 8125 27285 8159 27319
rect 9045 27285 9079 27319
rect 11253 27285 11287 27319
rect 13093 27285 13127 27319
rect 13369 27285 13403 27319
rect 13461 27285 13495 27319
rect 15025 27285 15059 27319
rect 19441 27285 19475 27319
rect 19901 27285 19935 27319
rect 20085 27285 20119 27319
rect 21925 27285 21959 27319
rect 25605 27285 25639 27319
rect 29377 27285 29411 27319
rect 6377 27081 6411 27115
rect 6545 27081 6579 27115
rect 7021 27081 7055 27115
rect 9597 27081 9631 27115
rect 12449 27081 12483 27115
rect 14013 27081 14047 27115
rect 21281 27081 21315 27115
rect 22661 27081 22695 27115
rect 27721 27081 27755 27115
rect 28917 27081 28951 27115
rect 6745 27013 6779 27047
rect 8125 27013 8159 27047
rect 29285 27013 29319 27047
rect 6929 26945 6963 26979
rect 7113 26945 7147 26979
rect 7849 26945 7883 26979
rect 9781 26945 9815 26979
rect 12357 26945 12391 26979
rect 13277 26945 13311 26979
rect 14105 26945 14139 26979
rect 14841 26945 14875 26979
rect 15209 26945 15243 26979
rect 18521 26945 18555 26979
rect 18705 26945 18739 26979
rect 21189 26945 21223 26979
rect 22569 26945 22603 26979
rect 25237 26945 25271 26979
rect 27353 26945 27387 26979
rect 29009 26945 29043 26979
rect 9873 26877 9907 26911
rect 13369 26877 13403 26911
rect 24961 26877 24995 26911
rect 27445 26877 27479 26911
rect 6561 26741 6595 26775
rect 15209 26741 15243 26775
rect 15393 26741 15427 26775
rect 18521 26741 18555 26775
rect 23489 26741 23523 26775
rect 29193 26741 29227 26775
rect 18061 26537 18095 26571
rect 20269 26537 20303 26571
rect 20545 26537 20579 26571
rect 23765 26537 23799 26571
rect 24041 26537 24075 26571
rect 29193 26537 29227 26571
rect 11161 26469 11195 26503
rect 16037 26469 16071 26503
rect 20729 26469 20763 26503
rect 23489 26469 23523 26503
rect 27445 26469 27479 26503
rect 27997 26469 28031 26503
rect 11805 26401 11839 26435
rect 13185 26401 13219 26435
rect 14657 26401 14691 26435
rect 17233 26401 17267 26435
rect 18245 26401 18279 26435
rect 19349 26401 19383 26435
rect 24961 26401 24995 26435
rect 26709 26401 26743 26435
rect 27261 26401 27295 26435
rect 4261 26333 4295 26367
rect 4721 26333 4755 26367
rect 6469 26333 6503 26367
rect 6745 26333 6779 26367
rect 8401 26333 8435 26367
rect 9413 26333 9447 26367
rect 9505 26333 9539 26367
rect 10149 26333 10183 26367
rect 10333 26333 10367 26367
rect 10517 26333 10551 26367
rect 11345 26333 11379 26367
rect 11437 26333 11471 26367
rect 12633 26333 12667 26367
rect 12725 26333 12759 26367
rect 12909 26333 12943 26367
rect 13001 26333 13035 26367
rect 13093 26333 13127 26367
rect 13369 26333 13403 26367
rect 13461 26333 13495 26367
rect 15117 26333 15151 26367
rect 15301 26333 15335 26367
rect 15669 26333 15703 26367
rect 15853 26333 15887 26367
rect 16313 26333 16347 26367
rect 16957 26333 16991 26367
rect 17049 26333 17083 26367
rect 17325 26333 17359 26367
rect 17417 26333 17451 26367
rect 17510 26333 17544 26367
rect 17923 26333 17957 26367
rect 18337 26333 18371 26367
rect 18613 26333 18647 26367
rect 18705 26333 18739 26367
rect 18981 26333 19015 26367
rect 19257 26333 19291 26367
rect 19625 26333 19659 26367
rect 19809 26333 19843 26367
rect 20085 26333 20119 26367
rect 23213 26333 23247 26367
rect 23305 26333 23339 26367
rect 24041 26333 24075 26367
rect 24225 26333 24259 26367
rect 26985 26333 27019 26367
rect 27077 26333 27111 26367
rect 27169 26333 27203 26367
rect 27629 26333 27663 26367
rect 27721 26333 27755 26367
rect 1501 26265 1535 26299
rect 1685 26265 1719 26299
rect 4445 26265 4479 26299
rect 5825 26265 5859 26299
rect 6009 26265 6043 26299
rect 10609 26265 10643 26299
rect 10793 26265 10827 26299
rect 11713 26265 11747 26299
rect 16037 26265 16071 26299
rect 16221 26265 16255 26299
rect 16773 26265 16807 26299
rect 17693 26265 17727 26299
rect 17785 26265 17819 26299
rect 18797 26265 18831 26299
rect 19901 26265 19935 26299
rect 20361 26265 20395 26299
rect 23489 26265 23523 26299
rect 23581 26265 23615 26299
rect 23781 26265 23815 26299
rect 25237 26265 25271 26299
rect 29285 26265 29319 26299
rect 4629 26197 4663 26231
rect 4813 26197 4847 26231
rect 6193 26197 6227 26231
rect 6377 26197 6411 26231
rect 6653 26197 6687 26231
rect 8309 26197 8343 26231
rect 9689 26197 9723 26231
rect 10977 26197 11011 26231
rect 12449 26197 12483 26231
rect 13645 26197 13679 26231
rect 18429 26197 18463 26231
rect 19809 26197 19843 26231
rect 20561 26197 20595 26231
rect 23949 26197 23983 26231
rect 26801 26197 26835 26231
rect 27813 26197 27847 26231
rect 5457 25993 5491 26027
rect 6193 25993 6227 26027
rect 10241 25993 10275 26027
rect 13553 25993 13587 26027
rect 14381 25993 14415 26027
rect 15209 25993 15243 26027
rect 15945 25993 15979 26027
rect 17877 25993 17911 26027
rect 21649 25993 21683 26027
rect 21833 25993 21867 26027
rect 24777 25993 24811 26027
rect 25513 25993 25547 26027
rect 26157 25993 26191 26027
rect 29377 25993 29411 26027
rect 5825 25925 5859 25959
rect 16681 25925 16715 25959
rect 17049 25925 17083 25959
rect 23305 25925 23339 25959
rect 25973 25925 26007 25959
rect 27353 25925 27387 25959
rect 3709 25857 3743 25891
rect 5641 25857 5675 25891
rect 5917 25857 5951 25891
rect 6009 25857 6043 25891
rect 6469 25857 6503 25891
rect 6653 25857 6687 25891
rect 7021 25857 7055 25891
rect 7573 25857 7607 25891
rect 7721 25857 7755 25891
rect 7849 25857 7883 25891
rect 7941 25857 7975 25891
rect 8079 25857 8113 25891
rect 8401 25857 8435 25891
rect 8493 25857 8527 25891
rect 8953 25857 8987 25891
rect 9229 25857 9263 25891
rect 9321 25857 9355 25891
rect 9505 25857 9539 25891
rect 9597 25857 9631 25891
rect 9873 25857 9907 25891
rect 10425 25857 10459 25891
rect 10793 25857 10827 25891
rect 10977 25857 11011 25891
rect 11529 25857 11563 25891
rect 11805 25857 11839 25891
rect 11989 25857 12023 25891
rect 12265 25857 12299 25891
rect 12449 25857 12483 25891
rect 12817 25857 12851 25891
rect 13277 25857 13311 25891
rect 13369 25857 13403 25891
rect 13645 25857 13679 25891
rect 14105 25857 14139 25891
rect 14565 25857 14599 25891
rect 14749 25857 14783 25891
rect 14933 25857 14967 25891
rect 15117 25857 15151 25891
rect 15393 25857 15427 25891
rect 15485 25857 15519 25891
rect 15669 25857 15703 25891
rect 15761 25857 15795 25891
rect 16129 25857 16163 25891
rect 16497 25857 16531 25891
rect 16865 25857 16899 25891
rect 17141 25857 17175 25891
rect 18061 25857 18095 25891
rect 18153 25857 18187 25891
rect 18429 25857 18463 25891
rect 18521 25857 18555 25891
rect 19257 25857 19291 25891
rect 19349 25857 19383 25891
rect 19717 25857 19751 25891
rect 19809 25857 19843 25891
rect 19901 25857 19935 25891
rect 23581 25857 23615 25891
rect 24869 25857 24903 25891
rect 26249 25857 26283 25891
rect 27169 25857 27203 25891
rect 3985 25789 4019 25823
rect 6745 25789 6779 25823
rect 6837 25789 6871 25823
rect 9045 25789 9079 25823
rect 10609 25789 10643 25823
rect 10701 25789 10735 25823
rect 13001 25789 13035 25823
rect 13093 25789 13127 25823
rect 14841 25789 14875 25823
rect 18613 25789 18647 25823
rect 19533 25789 19567 25823
rect 20177 25789 20211 25823
rect 27629 25789 27663 25823
rect 27905 25789 27939 25823
rect 8217 25721 8251 25755
rect 10149 25721 10183 25755
rect 12357 25721 12391 25755
rect 12909 25721 12943 25755
rect 13369 25721 13403 25755
rect 18337 25721 18371 25755
rect 19165 25721 19199 25755
rect 25697 25721 25731 25755
rect 7205 25653 7239 25687
rect 9965 25653 9999 25687
rect 11989 25653 12023 25687
rect 12173 25653 12207 25687
rect 12633 25653 12667 25687
rect 14197 25653 14231 25687
rect 16405 25653 16439 25687
rect 27537 25653 27571 25687
rect 4169 25449 4203 25483
rect 4353 25449 4387 25483
rect 9965 25449 9999 25483
rect 11897 25449 11931 25483
rect 12909 25449 12943 25483
rect 14473 25449 14507 25483
rect 16313 25449 16347 25483
rect 17601 25449 17635 25483
rect 18521 25449 18555 25483
rect 21465 25449 21499 25483
rect 22293 25449 22327 25483
rect 27353 25449 27387 25483
rect 27997 25449 28031 25483
rect 28825 25449 28859 25483
rect 7849 25381 7883 25415
rect 11345 25381 11379 25415
rect 13553 25381 13587 25415
rect 7113 25313 7147 25347
rect 10885 25313 10919 25347
rect 14657 25313 14691 25347
rect 15945 25313 15979 25347
rect 17141 25313 17175 25347
rect 17233 25313 17267 25347
rect 27629 25313 27663 25347
rect 4721 25245 4755 25279
rect 6193 25245 6227 25279
rect 6341 25245 6375 25279
rect 6699 25245 6733 25279
rect 7021 25245 7055 25279
rect 7205 25245 7239 25279
rect 7573 25245 7607 25279
rect 7665 25245 7699 25279
rect 7941 25245 7975 25279
rect 8677 25245 8711 25279
rect 9413 25245 9447 25279
rect 9689 25245 9723 25279
rect 9781 25245 9815 25279
rect 10793 25245 10827 25279
rect 11069 25245 11103 25279
rect 11161 25245 11195 25279
rect 11437 25245 11471 25279
rect 11713 25245 11747 25279
rect 13093 25245 13127 25279
rect 13461 25245 13495 25279
rect 13553 25245 13587 25279
rect 13737 25245 13771 25279
rect 14565 25245 14599 25279
rect 15853 25245 15887 25279
rect 16129 25245 16163 25279
rect 16865 25245 16899 25279
rect 17049 25245 17083 25279
rect 17417 25245 17451 25279
rect 18613 25245 18647 25279
rect 19901 25245 19935 25279
rect 21557 25245 21591 25279
rect 22201 25245 22235 25279
rect 23397 25245 23431 25279
rect 23673 25245 23707 25279
rect 27261 25245 27295 25279
rect 27445 25245 27479 25279
rect 27813 25245 27847 25279
rect 28917 25245 28951 25279
rect 6469 25177 6503 25211
rect 6561 25177 6595 25211
rect 9597 25177 9631 25211
rect 13185 25177 13219 25211
rect 13277 25177 13311 25211
rect 14197 25177 14231 25211
rect 4353 25109 4387 25143
rect 6837 25109 6871 25143
rect 7389 25109 7423 25143
rect 8585 25109 8619 25143
rect 11529 25109 11563 25143
rect 14289 25109 14323 25143
rect 19809 25109 19843 25143
rect 23213 25109 23247 25143
rect 23581 25109 23615 25143
rect 5641 24905 5675 24939
rect 6653 24905 6687 24939
rect 15761 24905 15795 24939
rect 16681 24905 16715 24939
rect 17417 24905 17451 24939
rect 24133 24905 24167 24939
rect 7757 24837 7791 24871
rect 23825 24837 23859 24871
rect 24041 24837 24075 24871
rect 27353 24837 27387 24871
rect 1409 24769 1443 24803
rect 5582 24769 5616 24803
rect 6101 24769 6135 24803
rect 6837 24769 6871 24803
rect 7113 24769 7147 24803
rect 7941 24769 7975 24803
rect 10057 24769 10091 24803
rect 14657 24769 14691 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 15485 24769 15519 24803
rect 15577 24769 15611 24803
rect 16865 24769 16899 24803
rect 16957 24769 16991 24803
rect 17233 24769 17267 24803
rect 17325 24769 17359 24803
rect 17509 24769 17543 24803
rect 17601 24769 17635 24803
rect 18705 24769 18739 24803
rect 18889 24769 18923 24803
rect 18981 24769 19015 24803
rect 19073 24769 19107 24803
rect 19809 24769 19843 24803
rect 21833 24769 21867 24803
rect 26249 24769 26283 24803
rect 27261 24769 27295 24803
rect 27445 24769 27479 24803
rect 29285 24769 29319 24803
rect 7021 24701 7055 24735
rect 22109 24701 22143 24735
rect 23581 24701 23615 24735
rect 25605 24701 25639 24735
rect 25881 24701 25915 24735
rect 5457 24633 5491 24667
rect 19901 24633 19935 24667
rect 27629 24633 27663 24667
rect 1593 24565 1627 24599
rect 6009 24565 6043 24599
rect 6929 24565 6963 24599
rect 8125 24565 8159 24599
rect 9965 24565 9999 24599
rect 14749 24565 14783 24599
rect 17141 24565 17175 24599
rect 17693 24565 17727 24599
rect 19257 24565 19291 24599
rect 23673 24565 23707 24599
rect 23857 24565 23891 24599
rect 26341 24565 26375 24599
rect 27077 24565 27111 24599
rect 29193 24565 29227 24599
rect 2132 24361 2166 24395
rect 3985 24361 4019 24395
rect 4169 24361 4203 24395
rect 4997 24361 5031 24395
rect 5365 24361 5399 24395
rect 7573 24361 7607 24395
rect 17417 24361 17451 24395
rect 22477 24361 22511 24395
rect 22937 24361 22971 24395
rect 24225 24361 24259 24395
rect 25237 24361 25271 24395
rect 27169 24361 27203 24395
rect 4537 24293 4571 24327
rect 8677 24293 8711 24327
rect 9597 24293 9631 24327
rect 14749 24293 14783 24327
rect 15761 24293 15795 24327
rect 23121 24293 23155 24327
rect 1869 24225 1903 24259
rect 14105 24225 14139 24259
rect 14197 24225 14231 24259
rect 18797 24225 18831 24259
rect 19809 24225 19843 24259
rect 20453 24225 20487 24259
rect 21649 24225 21683 24259
rect 22109 24225 22143 24259
rect 23765 24225 23799 24259
rect 25421 24225 25455 24259
rect 4813 24157 4847 24191
rect 4905 24157 4939 24191
rect 5089 24157 5123 24191
rect 5273 24157 5307 24191
rect 5457 24157 5491 24191
rect 5917 24157 5951 24191
rect 6065 24157 6099 24191
rect 6285 24157 6319 24191
rect 6382 24157 6416 24191
rect 7757 24157 7791 24191
rect 7849 24157 7883 24191
rect 8125 24157 8159 24191
rect 8401 24157 8435 24191
rect 8553 24157 8587 24191
rect 8769 24157 8803 24191
rect 8953 24157 8987 24191
rect 9137 24157 9171 24191
rect 9229 24157 9263 24191
rect 9321 24157 9355 24191
rect 9689 24157 9723 24191
rect 9873 24157 9907 24191
rect 9965 24157 9999 24191
rect 10057 24157 10091 24191
rect 10333 24157 10367 24191
rect 10701 24157 10735 24191
rect 11897 24157 11931 24191
rect 11990 24157 12024 24191
rect 12173 24157 12207 24191
rect 12265 24157 12299 24191
rect 12362 24157 12396 24191
rect 12817 24157 12851 24191
rect 13185 24157 13219 24191
rect 14568 24157 14602 24191
rect 15025 24157 15059 24191
rect 15301 24157 15335 24191
rect 15393 24157 15427 24191
rect 15669 24157 15703 24191
rect 15853 24157 15887 24191
rect 16865 24157 16899 24191
rect 16957 24157 16991 24191
rect 17213 24157 17247 24191
rect 17509 24157 17543 24191
rect 18061 24157 18095 24191
rect 18429 24157 18463 24191
rect 18521 24157 18555 24191
rect 18889 24157 18923 24191
rect 19625 24157 19659 24191
rect 19901 24157 19935 24191
rect 19993 24157 20027 24191
rect 20177 24157 20211 24191
rect 20545 24157 20579 24191
rect 21005 24157 21039 24191
rect 21373 24157 21407 24191
rect 21833 24157 21867 24191
rect 21925 24157 21959 24191
rect 22201 24157 22235 24191
rect 22385 24157 22419 24191
rect 23857 24157 23891 24191
rect 25329 24157 25363 24191
rect 27629 24157 27663 24191
rect 4721 24089 4755 24123
rect 6193 24089 6227 24123
rect 7941 24089 7975 24123
rect 8217 24089 8251 24123
rect 10517 24089 10551 24123
rect 10609 24089 10643 24123
rect 12909 24089 12943 24123
rect 13001 24089 13035 24123
rect 15209 24089 15243 24123
rect 17049 24089 17083 24123
rect 17969 24089 18003 24123
rect 21189 24089 21223 24123
rect 21281 24089 21315 24123
rect 23397 24089 23431 24123
rect 25697 24089 25731 24123
rect 27905 24089 27939 24123
rect 3617 24021 3651 24055
rect 4169 24021 4203 24055
rect 6561 24021 6595 24055
rect 10241 24021 10275 24055
rect 10885 24021 10919 24055
rect 12541 24021 12575 24055
rect 12633 24021 12667 24055
rect 14565 24021 14599 24055
rect 15577 24021 15611 24055
rect 16681 24021 16715 24055
rect 18153 24021 18187 24055
rect 18613 24021 18647 24055
rect 19441 24021 19475 24055
rect 20269 24021 20303 24055
rect 20913 24021 20947 24055
rect 21557 24021 21591 24055
rect 29377 24021 29411 24055
rect 3249 23817 3283 23851
rect 4261 23817 4295 23851
rect 4629 23817 4663 23851
rect 7757 23817 7791 23851
rect 9873 23817 9907 23851
rect 11345 23817 11379 23851
rect 13277 23817 13311 23851
rect 14473 23817 14507 23851
rect 19717 23817 19751 23851
rect 26341 23817 26375 23851
rect 28181 23817 28215 23851
rect 28917 23817 28951 23851
rect 4997 23749 5031 23783
rect 8861 23749 8895 23783
rect 11161 23749 11195 23783
rect 12725 23749 12759 23783
rect 14105 23749 14139 23783
rect 14197 23749 14231 23783
rect 16865 23749 16899 23783
rect 18429 23749 18463 23783
rect 19901 23749 19935 23783
rect 29101 23749 29135 23783
rect 29285 23749 29319 23783
rect 1409 23681 1443 23715
rect 3341 23681 3375 23715
rect 4169 23681 4203 23715
rect 4353 23681 4387 23715
rect 4721 23681 4755 23715
rect 4813 23681 4847 23715
rect 5917 23681 5951 23715
rect 6653 23681 6687 23715
rect 7021 23681 7055 23715
rect 7205 23681 7239 23715
rect 7297 23681 7331 23715
rect 7389 23681 7423 23715
rect 7665 23681 7699 23715
rect 8309 23681 8343 23715
rect 8585 23681 8619 23715
rect 8677 23681 8711 23715
rect 9321 23681 9355 23715
rect 9505 23681 9539 23715
rect 9597 23681 9631 23715
rect 9689 23681 9723 23715
rect 9965 23681 9999 23715
rect 10057 23681 10091 23715
rect 10241 23681 10275 23715
rect 10517 23681 10551 23715
rect 10701 23681 10735 23715
rect 10793 23681 10827 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 11989 23681 12023 23715
rect 12173 23681 12207 23715
rect 13001 23681 13035 23715
rect 13093 23681 13127 23715
rect 13369 23681 13403 23715
rect 13829 23681 13863 23715
rect 13922 23681 13956 23715
rect 14335 23681 14369 23715
rect 17049 23681 17083 23715
rect 18889 23681 18923 23715
rect 19625 23681 19659 23715
rect 20269 23681 20303 23715
rect 20637 23681 20671 23715
rect 26801 23681 26835 23715
rect 27169 23681 27203 23715
rect 27445 23681 27479 23715
rect 27813 23681 27847 23715
rect 29009 23681 29043 23715
rect 1685 23613 1719 23647
rect 10425 23613 10459 23647
rect 12633 23613 12667 23647
rect 18797 23613 18831 23647
rect 27261 23613 27295 23647
rect 27353 23613 27387 23647
rect 27721 23613 27755 23647
rect 7573 23545 7607 23579
rect 8401 23545 8435 23579
rect 20085 23545 20119 23579
rect 26525 23545 26559 23579
rect 26985 23545 27019 23579
rect 4445 23477 4479 23511
rect 6009 23477 6043 23511
rect 6745 23477 6779 23511
rect 10517 23477 10551 23511
rect 11161 23477 11195 23511
rect 13461 23477 13495 23511
rect 16681 23477 16715 23511
rect 18521 23477 18555 23511
rect 19073 23477 19107 23511
rect 19901 23477 19935 23511
rect 20545 23477 20579 23511
rect 4445 23273 4479 23307
rect 5917 23273 5951 23307
rect 8033 23273 8067 23307
rect 12265 23273 12299 23307
rect 12909 23273 12943 23307
rect 15577 23273 15611 23307
rect 16129 23273 16163 23307
rect 16589 23273 16623 23307
rect 18981 23273 19015 23307
rect 21741 23273 21775 23307
rect 27261 23273 27295 23307
rect 8217 23205 8251 23239
rect 12725 23205 12759 23239
rect 15025 23205 15059 23239
rect 15853 23205 15887 23239
rect 17049 23205 17083 23239
rect 17325 23205 17359 23239
rect 12449 23137 12483 23171
rect 14381 23137 14415 23171
rect 15669 23137 15703 23171
rect 24685 23137 24719 23171
rect 24869 23137 24903 23171
rect 28273 23137 28307 23171
rect 4353 23069 4387 23103
rect 4537 23069 4571 23103
rect 5365 23069 5399 23103
rect 5733 23069 5767 23103
rect 7389 23069 7423 23103
rect 7482 23069 7516 23103
rect 7895 23069 7929 23103
rect 8309 23069 8343 23103
rect 10977 23069 11011 23103
rect 11069 23069 11103 23103
rect 11161 23069 11195 23103
rect 12541 23069 12575 23103
rect 12817 23069 12851 23103
rect 14105 23069 14139 23103
rect 14197 23069 14231 23103
rect 14473 23069 14507 23103
rect 14841 23069 14875 23103
rect 15301 23069 15335 23103
rect 15393 23069 15427 23103
rect 15945 23069 15979 23103
rect 16405 23069 16439 23103
rect 16681 23071 16715 23105
rect 16773 23069 16807 23103
rect 17141 23069 17175 23103
rect 17325 23069 17359 23103
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 18061 23069 18095 23103
rect 18153 23069 18187 23103
rect 18705 23069 18739 23103
rect 18797 23069 18831 23103
rect 19073 23069 19107 23103
rect 21281 23069 21315 23103
rect 24501 23069 24535 23103
rect 24593 23069 24627 23103
rect 25145 23069 25179 23103
rect 27169 23069 27203 23103
rect 27353 23069 27387 23103
rect 27813 23069 27847 23103
rect 28089 23069 28123 23103
rect 5549 23001 5583 23035
rect 5641 23001 5675 23035
rect 7665 23001 7699 23035
rect 7757 23001 7791 23035
rect 11345 23001 11379 23035
rect 12265 23001 12299 23035
rect 14657 23001 14691 23035
rect 14749 23001 14783 23035
rect 15577 23001 15611 23035
rect 15669 23001 15703 23035
rect 16865 23001 16899 23035
rect 17049 23001 17083 23035
rect 18521 23001 18555 23035
rect 23213 23001 23247 23035
rect 27445 23001 27479 23035
rect 27629 23001 27663 23035
rect 14381 22933 14415 22967
rect 15117 22933 15151 22967
rect 18429 22933 18463 22967
rect 25053 22933 25087 22967
rect 27905 22933 27939 22967
rect 4537 22729 4571 22763
rect 9045 22729 9079 22763
rect 9873 22729 9907 22763
rect 16681 22729 16715 22763
rect 18981 22729 19015 22763
rect 21189 22729 21223 22763
rect 25421 22729 25455 22763
rect 29377 22729 29411 22763
rect 5089 22661 5123 22695
rect 5549 22661 5583 22695
rect 6101 22661 6135 22695
rect 7665 22661 7699 22695
rect 10517 22661 10551 22695
rect 13001 22661 13035 22695
rect 17233 22661 17267 22695
rect 17325 22661 17359 22695
rect 17877 22661 17911 22695
rect 17969 22661 18003 22695
rect 18337 22661 18371 22695
rect 19257 22661 19291 22695
rect 21557 22661 21591 22695
rect 23949 22661 23983 22695
rect 27905 22661 27939 22695
rect 1685 22593 1719 22627
rect 2789 22593 2823 22627
rect 4905 22593 4939 22627
rect 5365 22593 5399 22627
rect 5641 22593 5675 22627
rect 5733 22593 5767 22627
rect 6193 22593 6227 22627
rect 6377 22593 6411 22627
rect 7549 22593 7583 22627
rect 7757 22593 7791 22627
rect 7895 22593 7929 22627
rect 9137 22593 9171 22627
rect 9965 22593 9999 22627
rect 10609 22593 10643 22627
rect 10793 22593 10827 22627
rect 10977 22593 11011 22627
rect 11621 22593 11655 22627
rect 12817 22593 12851 22627
rect 12909 22593 12943 22627
rect 13185 22593 13219 22627
rect 16957 22593 16991 22627
rect 17601 22593 17635 22627
rect 17694 22593 17728 22627
rect 18107 22593 18141 22627
rect 18521 22593 18555 22627
rect 18613 22593 18647 22627
rect 18889 22593 18923 22627
rect 19165 22593 19199 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 19809 22593 19843 22627
rect 19993 22593 20027 22627
rect 20361 22593 20395 22627
rect 20637 22593 20671 22627
rect 20913 22593 20947 22627
rect 21005 22593 21039 22627
rect 21465 22593 21499 22627
rect 21833 22593 21867 22627
rect 23673 22593 23707 22627
rect 27169 22593 27203 22627
rect 1409 22525 1443 22559
rect 3065 22525 3099 22559
rect 6469 22525 6503 22559
rect 16865 22525 16899 22559
rect 18797 22525 18831 22559
rect 20085 22525 20119 22559
rect 20177 22525 20211 22559
rect 22109 22525 22143 22559
rect 27629 22525 27663 22559
rect 18245 22457 18279 22491
rect 4721 22389 4755 22423
rect 5917 22389 5951 22423
rect 7389 22389 7423 22423
rect 10977 22389 11011 22423
rect 11713 22389 11747 22423
rect 12633 22389 12667 22423
rect 20545 22389 20579 22423
rect 20729 22389 20763 22423
rect 23581 22389 23615 22423
rect 27077 22389 27111 22423
rect 4261 22185 4295 22219
rect 4445 22185 4479 22219
rect 14841 22185 14875 22219
rect 16957 22185 16991 22219
rect 20269 22185 20303 22219
rect 21170 22185 21204 22219
rect 24869 22185 24903 22219
rect 25310 22185 25344 22219
rect 27445 22185 27479 22219
rect 11345 22117 11379 22151
rect 14289 22117 14323 22151
rect 23305 22117 23339 22151
rect 3893 22049 3927 22083
rect 7665 22049 7699 22083
rect 7757 22049 7791 22083
rect 9229 22049 9263 22083
rect 9321 22049 9355 22083
rect 11529 22049 11563 22083
rect 12357 22049 12391 22083
rect 13369 22049 13403 22083
rect 14565 22049 14599 22083
rect 19533 22049 19567 22083
rect 20913 22049 20947 22083
rect 24501 22049 24535 22083
rect 25053 22049 25087 22083
rect 28917 22049 28951 22083
rect 3801 21981 3835 22015
rect 6193 21981 6227 22015
rect 6377 21981 6411 22015
rect 6469 21981 6503 22015
rect 6617 21981 6651 22015
rect 6745 21981 6779 22015
rect 6934 21981 6968 22015
rect 7389 21981 7423 22015
rect 7573 21981 7607 22015
rect 7941 21981 7975 22015
rect 8585 21981 8619 22015
rect 8953 21981 8987 22015
rect 9137 21981 9171 22015
rect 9505 21981 9539 22015
rect 9965 21981 9999 22015
rect 10057 21981 10091 22015
rect 10149 21981 10183 22015
rect 10333 21981 10367 22015
rect 10655 21981 10689 22015
rect 10793 21981 10827 22015
rect 11068 21981 11102 22015
rect 11161 21981 11195 22015
rect 11253 21981 11287 22015
rect 11800 21981 11834 22015
rect 12172 21981 12206 22015
rect 12265 21981 12299 22015
rect 12571 21981 12605 22015
rect 12725 21981 12759 22015
rect 13093 21981 13127 22015
rect 13185 21981 13219 22015
rect 13461 21981 13495 22015
rect 13553 21981 13587 22015
rect 13737 21981 13771 22015
rect 14197 21981 14231 22015
rect 14657 21981 14691 22015
rect 14749 21981 14783 22015
rect 15209 21981 15243 22015
rect 16865 21981 16899 22015
rect 19441 21981 19475 22015
rect 19717 21981 19751 22015
rect 20085 21981 20119 22015
rect 22937 21981 22971 22015
rect 24593 21981 24627 22015
rect 27077 21981 27111 22015
rect 27261 21981 27295 22015
rect 29009 21981 29043 22015
rect 29285 21981 29319 22015
rect 4629 21913 4663 21947
rect 6285 21913 6319 21947
rect 6837 21913 6871 21947
rect 8125 21913 8159 21947
rect 8217 21913 8251 21947
rect 8401 21913 8435 21947
rect 10885 21913 10919 21947
rect 11897 21913 11931 21947
rect 11989 21913 12023 21947
rect 13645 21913 13679 21947
rect 19901 21913 19935 21947
rect 19993 21913 20027 21947
rect 22845 21913 22879 21947
rect 23581 21913 23615 21947
rect 26893 21913 26927 21947
rect 4429 21845 4463 21879
rect 7113 21845 7147 21879
rect 9689 21845 9723 21879
rect 9781 21845 9815 21879
rect 10517 21845 10551 21879
rect 11529 21845 11563 21879
rect 11621 21845 11655 21879
rect 12909 21845 12943 21879
rect 15301 21845 15335 21879
rect 22661 21845 22695 21879
rect 23121 21845 23155 21879
rect 26801 21845 26835 21879
rect 27169 21845 27203 21879
rect 29193 21845 29227 21879
rect 8033 21641 8067 21675
rect 8585 21641 8619 21675
rect 9505 21641 9539 21675
rect 21189 21641 21223 21675
rect 21925 21641 21959 21675
rect 26433 21641 26467 21675
rect 29285 21641 29319 21675
rect 6745 21573 6779 21607
rect 7757 21573 7791 21607
rect 13185 21573 13219 21607
rect 14841 21573 14875 21607
rect 16313 21573 16347 21607
rect 16497 21573 16531 21607
rect 17417 21573 17451 21607
rect 18981 21573 19015 21607
rect 25421 21573 25455 21607
rect 1501 21505 1535 21539
rect 2881 21505 2915 21539
rect 5733 21505 5767 21539
rect 5917 21505 5951 21539
rect 6561 21505 6595 21539
rect 6653 21505 6687 21539
rect 6929 21505 6963 21539
rect 7481 21505 7515 21539
rect 7665 21505 7699 21539
rect 7849 21505 7883 21539
rect 8217 21505 8251 21539
rect 8401 21505 8435 21539
rect 8861 21505 8895 21539
rect 9413 21505 9447 21539
rect 9597 21505 9631 21539
rect 10701 21505 10735 21539
rect 11069 21505 11103 21539
rect 13001 21505 13035 21539
rect 13093 21505 13127 21539
rect 13369 21505 13403 21539
rect 14381 21505 14415 21539
rect 14565 21505 14599 21539
rect 14657 21505 14691 21539
rect 14933 21505 14967 21539
rect 15025 21505 15059 21539
rect 15301 21505 15335 21539
rect 16221 21505 16255 21539
rect 16865 21505 16899 21539
rect 16957 21505 16991 21539
rect 17233 21505 17267 21539
rect 17325 21505 17359 21539
rect 17509 21505 17543 21539
rect 18521 21505 18555 21539
rect 18797 21505 18831 21539
rect 19073 21505 19107 21539
rect 19165 21505 19199 21539
rect 21281 21505 21315 21539
rect 21833 21505 21867 21539
rect 22937 21505 22971 21539
rect 23121 21505 23155 21539
rect 23213 21505 23247 21539
rect 23357 21505 23391 21539
rect 23673 21505 23707 21539
rect 25513 21505 25547 21539
rect 25697 21505 25731 21539
rect 25881 21505 25915 21539
rect 26157 21505 26191 21539
rect 26249 21505 26283 21539
rect 26433 21505 26467 21539
rect 26617 21505 26651 21539
rect 26985 21505 27019 21539
rect 27537 21505 27571 21539
rect 3157 21437 3191 21471
rect 4905 21437 4939 21471
rect 10793 21437 10827 21471
rect 15393 21437 15427 21471
rect 15577 21437 15611 21471
rect 27445 21437 27479 21471
rect 27813 21437 27847 21471
rect 1685 21369 1719 21403
rect 5917 21369 5951 21403
rect 8769 21369 8803 21403
rect 10977 21369 11011 21403
rect 15209 21369 15243 21403
rect 16497 21369 16531 21403
rect 18613 21369 18647 21403
rect 27353 21369 27387 21403
rect 6377 21301 6411 21335
rect 8217 21301 8251 21335
rect 10609 21301 10643 21335
rect 11069 21301 11103 21335
rect 12817 21301 12851 21335
rect 14565 21301 14599 21335
rect 15485 21301 15519 21335
rect 16681 21301 16715 21335
rect 17141 21301 17175 21335
rect 19349 21301 19383 21335
rect 23489 21301 23523 21335
rect 25973 21301 26007 21335
rect 4077 21097 4111 21131
rect 9137 21097 9171 21131
rect 9965 21097 9999 21131
rect 12909 21097 12943 21131
rect 17969 21097 18003 21131
rect 23213 21097 23247 21131
rect 26801 21097 26835 21131
rect 27445 21097 27479 21131
rect 28733 21097 28767 21131
rect 12173 21029 12207 21063
rect 23581 21029 23615 21063
rect 19717 20961 19751 20995
rect 19809 20961 19843 20995
rect 20177 20961 20211 20995
rect 21465 20961 21499 20995
rect 23949 20961 23983 20995
rect 25053 20961 25087 20995
rect 27169 20961 27203 20995
rect 4169 20893 4203 20927
rect 6096 20893 6130 20927
rect 6468 20893 6502 20927
rect 6561 20893 6595 20927
rect 6837 20893 6871 20927
rect 9229 20893 9263 20927
rect 9321 20893 9355 20927
rect 9414 20893 9448 20927
rect 9827 20893 9861 20927
rect 10057 20893 10091 20927
rect 11897 20893 11931 20927
rect 12173 20893 12207 20927
rect 12817 20893 12851 20927
rect 16405 20893 16439 20927
rect 16589 20893 16623 20927
rect 16865 20893 16899 20927
rect 17049 20893 17083 20927
rect 17969 20893 18003 20927
rect 18061 20893 18095 20927
rect 19441 20893 19475 20927
rect 19625 20893 19659 20927
rect 19993 20893 20027 20927
rect 20448 20893 20482 20927
rect 20820 20893 20854 20927
rect 20913 20893 20947 20927
rect 21005 20893 21039 20927
rect 24409 20893 24443 20927
rect 24685 20893 24719 20927
rect 24777 20893 24811 20927
rect 26985 20893 27019 20927
rect 27077 20893 27111 20927
rect 27261 20893 27295 20927
rect 28825 20893 28859 20927
rect 29285 20893 29319 20927
rect 6193 20825 6227 20859
rect 6285 20825 6319 20859
rect 6929 20825 6963 20859
rect 8677 20825 8711 20859
rect 9597 20825 9631 20859
rect 9689 20825 9723 20859
rect 11805 20825 11839 20859
rect 18245 20825 18279 20859
rect 20545 20825 20579 20859
rect 20637 20825 20671 20859
rect 21189 20825 21223 20859
rect 21741 20825 21775 20859
rect 24593 20825 24627 20859
rect 25329 20825 25363 20859
rect 5917 20757 5951 20791
rect 6745 20757 6779 20791
rect 11989 20757 12023 20791
rect 16773 20757 16807 20791
rect 16865 20757 16899 20791
rect 17785 20757 17819 20791
rect 20269 20757 20303 20791
rect 21373 20757 21407 20791
rect 23489 20757 23523 20791
rect 24961 20757 24995 20791
rect 29193 20757 29227 20791
rect 9413 20553 9447 20587
rect 13001 20553 13035 20587
rect 13461 20553 13495 20587
rect 14289 20553 14323 20587
rect 15117 20553 15151 20587
rect 19073 20553 19107 20587
rect 21465 20553 21499 20587
rect 22569 20553 22603 20587
rect 24501 20553 24535 20587
rect 26157 20553 26191 20587
rect 7757 20485 7791 20519
rect 9045 20485 9079 20519
rect 9873 20485 9907 20519
rect 11805 20485 11839 20519
rect 13829 20485 13863 20519
rect 14749 20485 14783 20519
rect 14841 20485 14875 20519
rect 16037 20485 16071 20519
rect 23029 20485 23063 20519
rect 24685 20485 24719 20519
rect 3525 20417 3559 20451
rect 5641 20417 5675 20451
rect 5917 20417 5951 20451
rect 7021 20417 7055 20451
rect 8033 20417 8067 20451
rect 8309 20417 8343 20451
rect 8769 20417 8803 20451
rect 8917 20417 8951 20451
rect 9137 20417 9171 20451
rect 9234 20417 9268 20451
rect 9505 20417 9539 20451
rect 10977 20417 11011 20451
rect 11897 20417 11931 20451
rect 11989 20417 12023 20451
rect 12541 20417 12575 20451
rect 13093 20417 13127 20451
rect 13369 20417 13403 20451
rect 13461 20417 13495 20451
rect 13553 20417 13587 20451
rect 13737 20417 13771 20451
rect 13921 20417 13955 20451
rect 14197 20417 14231 20451
rect 14381 20417 14415 20451
rect 14473 20417 14507 20451
rect 14566 20417 14600 20451
rect 14938 20417 14972 20451
rect 15209 20417 15243 20451
rect 15393 20417 15427 20451
rect 16221 20417 16255 20451
rect 16313 20417 16347 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 17233 20417 17267 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 18245 20417 18279 20451
rect 18429 20417 18463 20451
rect 19257 20417 19291 20451
rect 19349 20417 19383 20451
rect 19534 20417 19568 20451
rect 19901 20417 19935 20451
rect 19993 20417 20027 20451
rect 20177 20417 20211 20451
rect 20269 20417 20303 20451
rect 20913 20417 20947 20451
rect 21097 20417 21131 20451
rect 21189 20417 21223 20451
rect 21281 20417 21315 20451
rect 22477 20417 22511 20451
rect 24777 20417 24811 20451
rect 26065 20417 26099 20451
rect 27537 20417 27571 20451
rect 3801 20349 3835 20383
rect 5549 20349 5583 20383
rect 7849 20349 7883 20383
rect 9597 20349 9631 20383
rect 9689 20349 9723 20383
rect 11529 20349 11563 20383
rect 11621 20349 11655 20383
rect 12265 20349 12299 20383
rect 12884 20349 12918 20383
rect 15301 20349 15335 20383
rect 16957 20349 16991 20383
rect 17049 20349 17083 20383
rect 18153 20349 18187 20383
rect 19441 20349 19475 20383
rect 22753 20349 22787 20383
rect 27629 20349 27663 20383
rect 8401 20281 8435 20315
rect 12725 20281 12759 20315
rect 16497 20281 16531 20315
rect 18613 20281 18647 20315
rect 6009 20213 6043 20247
rect 6193 20213 6227 20247
rect 7757 20213 7791 20247
rect 8217 20213 8251 20247
rect 9689 20213 9723 20247
rect 12449 20213 12483 20247
rect 16313 20213 16347 20247
rect 17417 20213 17451 20247
rect 19717 20213 19751 20247
rect 27813 20213 27847 20247
rect 4537 20009 4571 20043
rect 6193 20009 6227 20043
rect 9045 20009 9079 20043
rect 16865 20009 16899 20043
rect 18337 20009 18371 20043
rect 20637 20009 20671 20043
rect 26709 20009 26743 20043
rect 29377 20009 29411 20043
rect 5917 19941 5951 19975
rect 10057 19941 10091 19975
rect 15301 19941 15335 19975
rect 18429 19941 18463 19975
rect 19717 19941 19751 19975
rect 19809 19941 19843 19975
rect 2789 19873 2823 19907
rect 6653 19873 6687 19907
rect 7481 19873 7515 19907
rect 11437 19873 11471 19907
rect 11621 19873 11655 19907
rect 11713 19873 11747 19907
rect 11897 19873 11931 19907
rect 20177 19873 20211 19907
rect 21557 19873 21591 19907
rect 22109 19873 22143 19907
rect 24961 19873 24995 19907
rect 27169 19873 27203 19907
rect 27261 19873 27295 19907
rect 27629 19873 27663 19907
rect 27905 19873 27939 19907
rect 1501 19805 1535 19839
rect 1685 19805 1719 19839
rect 4445 19805 4479 19839
rect 5825 19805 5859 19839
rect 6285 19805 6319 19839
rect 6377 19805 6411 19839
rect 6561 19805 6595 19839
rect 6745 19805 6779 19839
rect 6929 19805 6963 19839
rect 7389 19805 7423 19839
rect 7665 19805 7699 19839
rect 7757 19805 7791 19839
rect 8217 19805 8251 19839
rect 8401 19805 8435 19839
rect 8585 19805 8619 19839
rect 8953 19805 8987 19839
rect 9965 19805 9999 19839
rect 10149 19805 10183 19839
rect 10241 19805 10275 19839
rect 10425 19805 10459 19839
rect 10701 19805 10735 19839
rect 10793 19805 10827 19839
rect 10977 19805 11011 19839
rect 11161 19805 11195 19839
rect 11805 19805 11839 19839
rect 12725 19805 12759 19839
rect 13001 19805 13035 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 14750 19805 14784 19839
rect 14933 19805 14967 19839
rect 15122 19805 15156 19839
rect 15577 19805 15611 19839
rect 16957 19805 16991 19839
rect 17693 19805 17727 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18613 19805 18647 19839
rect 18705 19805 18739 19839
rect 18981 19805 19015 19839
rect 19637 19805 19671 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 20361 19805 20395 19839
rect 20453 19805 20487 19839
rect 21097 19805 21131 19839
rect 21189 19805 21223 19839
rect 21833 19805 21867 19839
rect 21925 19805 21959 19839
rect 22201 19805 22235 19839
rect 26985 19805 27019 19839
rect 27077 19805 27111 19839
rect 2697 19737 2731 19771
rect 8309 19737 8343 19771
rect 11069 19737 11103 19771
rect 15025 19737 15059 19771
rect 15485 19737 15519 19771
rect 18797 19737 18831 19771
rect 19441 19737 19475 19771
rect 21465 19737 21499 19771
rect 25237 19737 25271 19771
rect 2237 19669 2271 19703
rect 2605 19669 2639 19703
rect 7113 19669 7147 19703
rect 7941 19669 7975 19703
rect 8033 19669 8067 19703
rect 10425 19669 10459 19703
rect 11345 19669 11379 19703
rect 12817 19669 12851 19703
rect 13185 19669 13219 19703
rect 14473 19669 14507 19703
rect 20913 19669 20947 19703
rect 21649 19669 21683 19703
rect 26801 19669 26835 19703
rect 7481 19465 7515 19499
rect 8769 19465 8803 19499
rect 9958 19465 9992 19499
rect 10885 19465 10919 19499
rect 12173 19465 12207 19499
rect 13001 19465 13035 19499
rect 18245 19465 18279 19499
rect 19809 19465 19843 19499
rect 20637 19465 20671 19499
rect 20827 19465 20861 19499
rect 20913 19465 20947 19499
rect 24685 19465 24719 19499
rect 25145 19465 25179 19499
rect 25973 19465 26007 19499
rect 27261 19465 27295 19499
rect 27353 19465 27387 19499
rect 27721 19465 27755 19499
rect 28917 19465 28951 19499
rect 1685 19397 1719 19431
rect 3433 19397 3467 19431
rect 5181 19397 5215 19431
rect 9873 19397 9907 19431
rect 11805 19397 11839 19431
rect 12633 19397 12667 19431
rect 17877 19397 17911 19431
rect 17969 19397 18003 19431
rect 19441 19397 19475 19431
rect 21373 19397 21407 19431
rect 24869 19397 24903 19431
rect 29285 19397 29319 19431
rect 1409 19329 1443 19363
rect 5089 19329 5123 19363
rect 6745 19329 6779 19363
rect 6929 19329 6963 19363
rect 7021 19329 7055 19363
rect 7297 19329 7331 19363
rect 8125 19329 8159 19363
rect 8309 19329 8343 19363
rect 8401 19329 8435 19363
rect 8493 19329 8527 19363
rect 8953 19329 8987 19363
rect 9321 19329 9355 19363
rect 9505 19329 9539 19363
rect 9781 19329 9815 19363
rect 10057 19329 10091 19363
rect 10793 19329 10827 19363
rect 10977 19329 11011 19363
rect 11897 19329 11931 19363
rect 12014 19329 12048 19363
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 12817 19329 12851 19363
rect 14289 19329 14323 19363
rect 14473 19329 14507 19363
rect 14841 19329 14875 19363
rect 16865 19329 16899 19363
rect 16957 19329 16991 19363
rect 17233 19329 17267 19363
rect 17693 19329 17727 19363
rect 18061 19329 18095 19363
rect 19257 19329 19291 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 19993 19329 20027 19363
rect 20086 19329 20120 19363
rect 20269 19329 20303 19363
rect 20361 19329 20395 19363
rect 20499 19329 20533 19363
rect 20729 19329 20763 19363
rect 21005 19329 21039 19363
rect 21465 19329 21499 19363
rect 22937 19329 22971 19363
rect 24961 19329 24995 19363
rect 25881 19329 25915 19363
rect 27169 19329 27203 19363
rect 27629 19329 27663 19363
rect 27813 19329 27847 19363
rect 29009 19329 29043 19363
rect 5273 19261 5307 19295
rect 7113 19261 7147 19295
rect 9229 19261 9263 19295
rect 11529 19261 11563 19295
rect 14565 19261 14599 19295
rect 14657 19261 14691 19295
rect 17141 19261 17175 19295
rect 23213 19261 23247 19295
rect 25605 19261 25639 19295
rect 26985 19261 27019 19295
rect 4721 19193 4755 19227
rect 9413 19193 9447 19227
rect 25329 19193 25363 19227
rect 27537 19193 27571 19227
rect 8677 19125 8711 19159
rect 9137 19125 9171 19159
rect 15025 19125 15059 19159
rect 16681 19125 16715 19159
rect 29193 19125 29227 19159
rect 2421 18921 2455 18955
rect 3801 18921 3835 18955
rect 6837 18921 6871 18955
rect 7205 18921 7239 18955
rect 7389 18921 7423 18955
rect 10517 18921 10551 18955
rect 18521 18921 18555 18955
rect 18613 18921 18647 18955
rect 21281 18921 21315 18955
rect 22477 18921 22511 18955
rect 5089 18853 5123 18887
rect 9597 18853 9631 18887
rect 10057 18853 10091 18887
rect 15301 18853 15335 18887
rect 1685 18785 1719 18819
rect 3985 18785 4019 18819
rect 4629 18785 4663 18819
rect 5181 18785 5215 18819
rect 5457 18785 5491 18819
rect 6837 18785 6871 18819
rect 8309 18785 8343 18819
rect 9045 18785 9079 18819
rect 10149 18785 10183 18819
rect 14197 18785 14231 18819
rect 17233 18785 17267 18819
rect 18521 18785 18555 18819
rect 22109 18785 22143 18819
rect 27721 18785 27755 18819
rect 29101 18785 29135 18819
rect 1409 18717 1443 18751
rect 2329 18717 2363 18751
rect 4077 18717 4111 18751
rect 4721 18717 4755 18751
rect 5549 18717 5583 18751
rect 7021 18717 7055 18751
rect 7297 18717 7331 18751
rect 8033 18717 8067 18751
rect 8125 18717 8159 18751
rect 8401 18717 8435 18751
rect 8953 18717 8987 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 9873 18717 9907 18751
rect 10333 18717 10367 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 14381 18717 14415 18751
rect 14473 18717 14507 18751
rect 14657 18717 14691 18751
rect 14749 18717 14783 18751
rect 15025 18717 15059 18751
rect 15117 18717 15151 18751
rect 15669 18717 15703 18751
rect 15853 18717 15887 18751
rect 17049 18717 17083 18751
rect 17325 18717 17359 18751
rect 17417 18717 17451 18751
rect 17601 18717 17635 18751
rect 17877 18717 17911 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 18705 18717 18739 18751
rect 20361 18717 20395 18751
rect 21373 18717 21407 18751
rect 22201 18717 22235 18751
rect 22753 18717 22787 18751
rect 22845 18717 22879 18751
rect 27813 18717 27847 18751
rect 27997 18717 28031 18751
rect 29377 18717 29411 18751
rect 4353 18649 4387 18683
rect 4445 18649 4479 18683
rect 6561 18649 6595 18683
rect 7849 18649 7883 18683
rect 15301 18649 15335 18683
rect 18337 18649 18371 18683
rect 27353 18649 27387 18683
rect 27537 18649 27571 18683
rect 14933 18581 14967 18615
rect 15853 18581 15887 18615
rect 16865 18581 16899 18615
rect 17693 18581 17727 18615
rect 20269 18581 20303 18615
rect 28181 18581 28215 18615
rect 2513 18377 2547 18411
rect 4077 18377 4111 18411
rect 13553 18377 13587 18411
rect 15393 18377 15427 18411
rect 17509 18377 17543 18411
rect 21005 18377 21039 18411
rect 25053 18377 25087 18411
rect 29377 18377 29411 18411
rect 1685 18309 1719 18343
rect 10793 18309 10827 18343
rect 13829 18309 13863 18343
rect 15184 18309 15218 18343
rect 16957 18309 16991 18343
rect 27905 18309 27939 18343
rect 1777 18241 1811 18275
rect 2145 18241 2179 18275
rect 3985 18241 4019 18275
rect 4261 18241 4295 18275
rect 10241 18241 10275 18275
rect 10977 18241 11011 18275
rect 11805 18241 11839 18275
rect 13921 18241 13955 18275
rect 16313 18241 16347 18275
rect 16681 18241 16715 18275
rect 16774 18241 16808 18275
rect 17049 18241 17083 18275
rect 17187 18241 17221 18275
rect 17693 18241 17727 18275
rect 17785 18241 17819 18275
rect 18061 18241 18095 18275
rect 18337 18241 18371 18275
rect 18429 18241 18463 18275
rect 18521 18241 18555 18275
rect 18705 18241 18739 18275
rect 21097 18241 21131 18275
rect 21373 18241 21407 18275
rect 21465 18241 21499 18275
rect 21649 18241 21683 18275
rect 21833 18241 21867 18275
rect 21925 18241 21959 18275
rect 22109 18241 22143 18275
rect 22201 18241 22235 18275
rect 22845 18241 22879 18275
rect 23305 18241 23339 18275
rect 25329 18241 25363 18275
rect 26249 18241 26283 18275
rect 27629 18241 27663 18275
rect 2237 18173 2271 18207
rect 10333 18173 10367 18207
rect 12081 18173 12115 18207
rect 15301 18173 15335 18207
rect 15669 18173 15703 18207
rect 16037 18173 16071 18207
rect 22385 18173 22419 18207
rect 22753 18173 22787 18207
rect 23581 18173 23615 18207
rect 25237 18173 25271 18207
rect 4261 18105 4295 18139
rect 15761 18105 15795 18139
rect 18153 18105 18187 18139
rect 21649 18105 21683 18139
rect 23213 18105 23247 18139
rect 10609 18037 10643 18071
rect 15025 18037 15059 18071
rect 16221 18037 16255 18071
rect 17325 18037 17359 18071
rect 17969 18037 18003 18071
rect 25605 18037 25639 18071
rect 26341 18037 26375 18071
rect 2329 17833 2363 17867
rect 3801 17833 3835 17867
rect 8125 17833 8159 17867
rect 10793 17833 10827 17867
rect 11805 17833 11839 17867
rect 16589 17833 16623 17867
rect 22109 17833 22143 17867
rect 24501 17833 24535 17867
rect 28825 17833 28859 17867
rect 2605 17765 2639 17799
rect 5181 17765 5215 17799
rect 8585 17765 8619 17799
rect 27445 17765 27479 17799
rect 3433 17697 3467 17731
rect 3985 17697 4019 17731
rect 4077 17697 4111 17731
rect 4813 17697 4847 17731
rect 5022 17697 5056 17731
rect 5733 17697 5767 17731
rect 8033 17697 8067 17731
rect 10701 17697 10735 17731
rect 12265 17697 12299 17731
rect 12357 17697 12391 17731
rect 16405 17697 16439 17731
rect 19257 17697 19291 17731
rect 21281 17697 21315 17731
rect 25237 17697 25271 17731
rect 2237 17629 2271 17663
rect 2421 17629 2455 17663
rect 2513 17629 2547 17663
rect 2690 17629 2724 17663
rect 2973 17629 3007 17663
rect 3341 17629 3375 17663
rect 3525 17629 3559 17663
rect 4169 17629 4203 17663
rect 4261 17629 4295 17663
rect 4537 17629 4571 17663
rect 5641 17629 5675 17663
rect 6009 17629 6043 17663
rect 8309 17629 8343 17663
rect 8401 17629 8435 17663
rect 8953 17629 8987 17663
rect 9137 17629 9171 17663
rect 10793 17629 10827 17663
rect 11253 17629 11287 17663
rect 15669 17629 15703 17663
rect 16681 17629 16715 17663
rect 21833 17629 21867 17663
rect 21925 17629 21959 17663
rect 24593 17629 24627 17663
rect 28917 17629 28951 17663
rect 2789 17561 2823 17595
rect 3157 17561 3191 17595
rect 4905 17561 4939 17595
rect 6285 17561 6319 17595
rect 8125 17561 8159 17595
rect 10517 17561 10551 17595
rect 11069 17561 11103 17595
rect 11437 17561 11471 17595
rect 15853 17561 15887 17595
rect 16405 17561 16439 17595
rect 21005 17561 21039 17595
rect 25513 17561 25547 17595
rect 27077 17561 27111 17595
rect 5273 17493 5307 17527
rect 9137 17493 9171 17527
rect 10977 17493 11011 17527
rect 12173 17493 12207 17527
rect 15485 17493 15519 17527
rect 26985 17493 27019 17527
rect 27537 17493 27571 17527
rect 3433 17289 3467 17323
rect 3988 17289 4022 17323
rect 4261 17289 4295 17323
rect 6929 17289 6963 17323
rect 7113 17289 7147 17323
rect 18613 17289 18647 17323
rect 19349 17289 19383 17323
rect 19717 17289 19751 17323
rect 20085 17289 20119 17323
rect 26525 17289 26559 17323
rect 29193 17289 29227 17323
rect 1501 17221 1535 17255
rect 7481 17221 7515 17255
rect 10333 17221 10367 17255
rect 11253 17221 11287 17255
rect 20545 17221 20579 17255
rect 21465 17221 21499 17255
rect 26433 17221 26467 17255
rect 26801 17221 26835 17255
rect 27721 17221 27755 17255
rect 3433 17153 3467 17187
rect 3617 17153 3651 17187
rect 3801 17153 3835 17187
rect 3893 17153 3927 17187
rect 4261 17153 4295 17187
rect 4445 17153 4479 17187
rect 4629 17153 4663 17187
rect 6837 17153 6871 17187
rect 7573 17153 7607 17187
rect 8309 17153 8343 17187
rect 9137 17153 9171 17187
rect 10241 17153 10275 17187
rect 10425 17153 10459 17187
rect 10563 17153 10597 17187
rect 10701 17153 10735 17187
rect 10793 17153 10827 17187
rect 10977 17153 11011 17187
rect 11345 17153 11379 17187
rect 12357 17153 12391 17187
rect 12541 17153 12575 17187
rect 12817 17153 12851 17187
rect 13093 17153 13127 17187
rect 13277 17153 13311 17187
rect 13461 17153 13495 17187
rect 14105 17153 14139 17187
rect 16221 17153 16255 17187
rect 18245 17153 18279 17187
rect 19993 17153 20027 17187
rect 20637 17153 20671 17187
rect 21649 17153 21683 17187
rect 21833 17153 21867 17187
rect 21926 17153 21960 17187
rect 22109 17153 22143 17187
rect 22201 17153 22235 17187
rect 22298 17153 22332 17187
rect 25605 17153 25639 17187
rect 25789 17153 25823 17187
rect 26249 17153 26283 17187
rect 26617 17153 26651 17187
rect 27445 17153 27479 17187
rect 1685 17085 1719 17119
rect 7665 17085 7699 17119
rect 8401 17085 8435 17119
rect 8769 17085 8803 17119
rect 9229 17085 9263 17119
rect 10057 17085 10091 17119
rect 10885 17085 10919 17119
rect 14013 17085 14047 17119
rect 18153 17085 18187 17119
rect 19165 17085 19199 17119
rect 19257 17085 19291 17119
rect 4123 17017 4157 17051
rect 4445 17017 4479 17051
rect 8677 17017 8711 17051
rect 13185 17017 13219 17051
rect 13001 16949 13035 16983
rect 16313 16949 16347 16983
rect 21281 16949 21315 16983
rect 22477 16949 22511 16983
rect 25421 16949 25455 16983
rect 1593 16745 1627 16779
rect 18153 16745 18187 16779
rect 20913 16745 20947 16779
rect 21189 16745 21223 16779
rect 21465 16745 21499 16779
rect 26893 16745 26927 16779
rect 27537 16745 27571 16779
rect 28641 16745 28675 16779
rect 22845 16677 22879 16711
rect 29101 16677 29135 16711
rect 7573 16609 7607 16643
rect 7849 16609 7883 16643
rect 15209 16609 15243 16643
rect 17233 16609 17267 16643
rect 20821 16609 20855 16643
rect 21557 16609 21591 16643
rect 22385 16609 22419 16643
rect 25145 16609 25179 16643
rect 27077 16609 27111 16643
rect 27169 16609 27203 16643
rect 27261 16609 27295 16643
rect 27353 16609 27387 16643
rect 1501 16541 1535 16575
rect 6561 16541 6595 16575
rect 7481 16541 7515 16575
rect 10241 16541 10275 16575
rect 10425 16541 10459 16575
rect 10609 16541 10643 16575
rect 10763 16541 10797 16575
rect 12725 16541 12759 16575
rect 12909 16541 12943 16575
rect 13093 16541 13127 16575
rect 14289 16541 14323 16575
rect 17417 16541 17451 16575
rect 17601 16541 17635 16575
rect 17687 16541 17721 16575
rect 17785 16541 17819 16575
rect 17969 16541 18003 16575
rect 18245 16541 18279 16575
rect 18429 16541 18463 16575
rect 21005 16541 21039 16575
rect 21649 16541 21683 16575
rect 21741 16541 21775 16575
rect 21925 16541 21959 16575
rect 22477 16541 22511 16575
rect 24225 16541 24259 16575
rect 24869 16541 24903 16575
rect 25053 16541 25087 16575
rect 28273 16541 28307 16575
rect 28733 16541 28767 16575
rect 29009 16541 29043 16575
rect 29285 16541 29319 16575
rect 13001 16473 13035 16507
rect 15485 16473 15519 16507
rect 20729 16473 20763 16507
rect 25421 16473 25455 16507
rect 6653 16405 6687 16439
rect 10333 16405 10367 16439
rect 10977 16405 11011 16439
rect 13277 16405 13311 16439
rect 14381 16405 14415 16439
rect 17509 16405 17543 16439
rect 18337 16405 18371 16439
rect 21281 16405 21315 16439
rect 21925 16405 21959 16439
rect 24133 16405 24167 16439
rect 25053 16405 25087 16439
rect 28457 16405 28491 16439
rect 28917 16405 28951 16439
rect 9229 16201 9263 16235
rect 10517 16201 10551 16235
rect 11345 16201 11379 16235
rect 12173 16201 12207 16235
rect 15577 16201 15611 16235
rect 16037 16201 16071 16235
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 20913 16201 20947 16235
rect 23029 16201 23063 16235
rect 25605 16201 25639 16235
rect 26249 16201 26283 16235
rect 29377 16201 29411 16235
rect 3709 16133 3743 16167
rect 4169 16133 4203 16167
rect 5549 16133 5583 16167
rect 8401 16133 8435 16167
rect 13553 16133 13587 16167
rect 15301 16133 15335 16167
rect 24501 16133 24535 16167
rect 1685 16065 1719 16099
rect 3985 16065 4019 16099
rect 4077 16065 4111 16099
rect 4353 16065 4387 16099
rect 4629 16065 4663 16099
rect 4813 16065 4847 16099
rect 5181 16065 5215 16099
rect 5273 16065 5307 16099
rect 5365 16065 5399 16099
rect 6377 16065 6411 16099
rect 8861 16065 8895 16099
rect 9137 16065 9171 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 9965 16065 9999 16099
rect 10057 16065 10091 16099
rect 10241 16065 10275 16099
rect 10341 16065 10375 16099
rect 10977 16065 11011 16099
rect 11713 16065 11747 16099
rect 12176 16065 12210 16099
rect 13277 16065 13311 16099
rect 15945 16065 15979 16099
rect 19165 16065 19199 16099
rect 19717 16065 19751 16099
rect 19993 16065 20027 16099
rect 20257 16065 20291 16099
rect 20361 16065 20395 16099
rect 20788 16065 20822 16099
rect 22385 16065 22419 16099
rect 25237 16065 25271 16099
rect 25421 16065 25455 16099
rect 26157 16065 26191 16099
rect 27169 16065 27203 16099
rect 1961 15997 1995 16031
rect 6653 15997 6687 16031
rect 8953 15997 8987 16031
rect 9597 15997 9631 16031
rect 10885 15997 10919 16031
rect 16129 15997 16163 16031
rect 18061 15997 18095 16031
rect 19073 15997 19107 16031
rect 19809 15997 19843 16031
rect 22109 15997 22143 16031
rect 24777 15997 24811 16031
rect 27261 15997 27295 16031
rect 27629 15997 27663 16031
rect 27905 15997 27939 16031
rect 3801 15929 3835 15963
rect 9413 15929 9447 15963
rect 17693 15929 17727 15963
rect 18797 15929 18831 15963
rect 21833 15929 21867 15963
rect 27537 15929 27571 15963
rect 4445 15861 4479 15895
rect 8493 15861 8527 15895
rect 9781 15861 9815 15895
rect 11805 15861 11839 15895
rect 12357 15861 12391 15895
rect 17601 15861 17635 15895
rect 19717 15861 19751 15895
rect 22109 15861 22143 15895
rect 1593 15657 1627 15691
rect 2605 15657 2639 15691
rect 3617 15657 3651 15691
rect 3893 15657 3927 15691
rect 5457 15657 5491 15691
rect 6561 15657 6595 15691
rect 9045 15657 9079 15691
rect 10517 15657 10551 15691
rect 11437 15657 11471 15691
rect 11805 15657 11839 15691
rect 13277 15657 13311 15691
rect 16681 15657 16715 15691
rect 18521 15657 18555 15691
rect 19717 15657 19751 15691
rect 19993 15657 20027 15691
rect 21005 15657 21039 15691
rect 4445 15589 4479 15623
rect 4813 15589 4847 15623
rect 13645 15589 13679 15623
rect 4721 15521 4755 15555
rect 7113 15521 7147 15555
rect 11529 15521 11563 15555
rect 17969 15521 18003 15555
rect 19349 15521 19383 15555
rect 20821 15521 20855 15555
rect 22109 15521 22143 15555
rect 23765 15521 23799 15555
rect 2513 15453 2547 15487
rect 3433 15453 3467 15487
rect 3617 15453 3651 15487
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 4353 15453 4387 15487
rect 4537 15453 4571 15487
rect 5273 15453 5307 15487
rect 5366 15453 5400 15487
rect 6929 15453 6963 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 10057 15453 10091 15487
rect 10333 15453 10367 15487
rect 11437 15453 11471 15487
rect 13001 15453 13035 15487
rect 13093 15453 13127 15487
rect 13461 15453 13495 15487
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 13921 15453 13955 15487
rect 14289 15453 14323 15487
rect 15025 15453 15059 15487
rect 15209 15453 15243 15487
rect 17325 15453 17359 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 17693 15453 17727 15487
rect 18061 15453 18095 15487
rect 18153 15453 18187 15487
rect 18337 15453 18371 15487
rect 18521 15453 18555 15487
rect 19441 15453 19475 15487
rect 19809 15453 19843 15487
rect 20729 15453 20763 15487
rect 21005 15453 21039 15487
rect 22201 15453 22235 15487
rect 23673 15453 23707 15487
rect 24593 15453 24627 15487
rect 27353 15453 27387 15487
rect 27537 15453 27571 15487
rect 29101 15453 29135 15487
rect 29377 15453 29411 15487
rect 1501 15385 1535 15419
rect 5181 15385 5215 15419
rect 7021 15385 7055 15419
rect 10149 15385 10183 15419
rect 15393 15385 15427 15419
rect 23581 15385 23615 15419
rect 12633 15317 12667 15351
rect 14381 15317 14415 15351
rect 21189 15317 21223 15351
rect 22569 15317 22603 15351
rect 23213 15317 23247 15351
rect 24501 15317 24535 15351
rect 27445 15317 27479 15351
rect 12725 15113 12759 15147
rect 13369 15113 13403 15147
rect 16957 15113 16991 15147
rect 27905 15113 27939 15147
rect 16313 15045 16347 15079
rect 23305 15045 23339 15079
rect 25053 15045 25087 15079
rect 27813 15045 27847 15079
rect 6653 14977 6687 15011
rect 6837 14977 6871 15011
rect 6929 14977 6963 15011
rect 7113 14977 7147 15011
rect 10149 14977 10183 15011
rect 11529 14977 11563 15011
rect 11713 14977 11747 15011
rect 11989 14977 12023 15011
rect 12357 14977 12391 15011
rect 12449 14977 12483 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 13277 14977 13311 15011
rect 13369 14977 13403 15011
rect 13553 14977 13587 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 17049 14977 17083 15011
rect 17233 14977 17267 15011
rect 22017 14977 22051 15011
rect 26157 14977 26191 15011
rect 27261 14977 27295 15011
rect 27997 14977 28031 15011
rect 28457 14977 28491 15011
rect 28549 14977 28583 15011
rect 14289 14909 14323 14943
rect 14565 14909 14599 14943
rect 21925 14909 21959 14943
rect 22385 14909 22419 14943
rect 23029 14909 23063 14943
rect 25881 14909 25915 14943
rect 27169 14909 27203 14943
rect 27353 14909 27387 14943
rect 27445 14909 27479 14943
rect 11897 14841 11931 14875
rect 13185 14841 13219 14875
rect 25605 14841 25639 14875
rect 26985 14841 27019 14875
rect 28181 14841 28215 14875
rect 6745 14773 6779 14807
rect 6929 14773 6963 14807
rect 10057 14773 10091 14807
rect 17233 14773 17267 14807
rect 25421 14773 25455 14807
rect 26065 14773 26099 14807
rect 27629 14773 27663 14807
rect 28273 14773 28307 14807
rect 6745 14569 6779 14603
rect 14289 14569 14323 14603
rect 15945 14569 15979 14603
rect 16221 14569 16255 14603
rect 26617 14569 26651 14603
rect 27537 14569 27571 14603
rect 27892 14569 27926 14603
rect 29377 14569 29411 14603
rect 6377 14501 6411 14535
rect 17969 14501 18003 14535
rect 18061 14501 18095 14535
rect 19349 14501 19383 14535
rect 4445 14433 4479 14467
rect 7021 14433 7055 14467
rect 8769 14433 8803 14467
rect 13461 14433 13495 14467
rect 15761 14433 15795 14467
rect 18337 14433 18371 14467
rect 18613 14433 18647 14467
rect 19073 14433 19107 14467
rect 24869 14433 24903 14467
rect 3433 14365 3467 14399
rect 9137 14365 9171 14399
rect 10057 14365 10091 14399
rect 10149 14365 10183 14399
rect 10425 14365 10459 14399
rect 10609 14365 10643 14399
rect 10977 14365 11011 14399
rect 13185 14365 13219 14399
rect 13277 14365 13311 14399
rect 13645 14365 13679 14399
rect 13829 14365 13863 14399
rect 14473 14365 14507 14399
rect 14657 14365 14691 14399
rect 14749 14365 14783 14399
rect 15669 14365 15703 14399
rect 16313 14365 16347 14399
rect 17509 14365 17543 14399
rect 17693 14365 17727 14399
rect 17877 14365 17911 14399
rect 18153 14365 18187 14399
rect 18705 14365 18739 14399
rect 19257 14365 19291 14399
rect 19441 14365 19475 14399
rect 19717 14365 19751 14399
rect 27629 14365 27663 14399
rect 4721 14297 4755 14331
rect 6745 14297 6779 14331
rect 7297 14297 7331 14331
rect 9045 14297 9079 14331
rect 10333 14297 10367 14331
rect 19993 14297 20027 14331
rect 21741 14297 21775 14331
rect 25145 14297 25179 14331
rect 27169 14297 27203 14331
rect 27353 14297 27387 14331
rect 3525 14229 3559 14263
rect 6193 14229 6227 14263
rect 6929 14229 6963 14263
rect 10517 14229 10551 14263
rect 10885 14229 10919 14263
rect 13461 14229 13495 14263
rect 13737 14229 13771 14263
rect 17601 14229 17635 14263
rect 5457 14025 5491 14059
rect 12173 14025 12207 14059
rect 12265 14025 12299 14059
rect 16037 14025 16071 14059
rect 16957 14025 16991 14059
rect 18337 14025 18371 14059
rect 18889 14025 18923 14059
rect 19809 14025 19843 14059
rect 20177 14025 20211 14059
rect 20269 14025 20303 14059
rect 20913 14025 20947 14059
rect 28917 14025 28951 14059
rect 4721 13957 4755 13991
rect 6561 13957 6595 13991
rect 6745 13957 6779 13991
rect 9413 13957 9447 13991
rect 9505 13957 9539 13991
rect 10885 13957 10919 13991
rect 12014 13957 12048 13991
rect 13093 13957 13127 13991
rect 14289 13957 14323 13991
rect 29101 13957 29135 13991
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 6837 13889 6871 13923
rect 7481 13889 7515 13923
rect 7573 13889 7607 13923
rect 9137 13889 9171 13923
rect 9229 13889 9263 13923
rect 9597 13889 9631 13923
rect 10609 13889 10643 13923
rect 10757 13889 10791 13923
rect 10977 13889 11011 13923
rect 11115 13889 11149 13923
rect 11529 13889 11563 13923
rect 12633 13889 12667 13923
rect 12955 13889 12989 13923
rect 13185 13889 13219 13923
rect 13368 13889 13402 13923
rect 13461 13889 13495 13923
rect 13737 13889 13771 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 14473 13889 14507 13923
rect 14657 13889 14691 13923
rect 16129 13889 16163 13923
rect 16865 13889 16899 13923
rect 17325 13889 17359 13923
rect 18245 13889 18279 13923
rect 18429 13889 18463 13923
rect 18521 13889 18555 13923
rect 18705 13889 18739 13923
rect 21005 13889 21039 13923
rect 22109 13889 22143 13923
rect 22569 13889 22603 13923
rect 29009 13889 29043 13923
rect 29285 13889 29319 13923
rect 1409 13821 1443 13855
rect 1685 13821 1719 13855
rect 2421 13821 2455 13855
rect 11805 13821 11839 13855
rect 11897 13821 11931 13855
rect 12541 13821 12575 13855
rect 13553 13821 13587 13855
rect 13921 13821 13955 13855
rect 14565 13821 14599 13855
rect 16221 13821 16255 13855
rect 17417 13821 17451 13855
rect 20361 13821 20395 13855
rect 22017 13821 22051 13855
rect 24593 13821 24627 13855
rect 24685 13821 24719 13855
rect 24961 13821 24995 13855
rect 27169 13821 27203 13855
rect 4537 13753 4571 13787
rect 6377 13753 6411 13787
rect 13829 13753 13863 13787
rect 27537 13753 27571 13787
rect 2684 13685 2718 13719
rect 4169 13685 4203 13719
rect 4721 13685 4755 13719
rect 6929 13685 6963 13719
rect 9045 13685 9079 13719
rect 9781 13685 9815 13719
rect 11253 13685 11287 13719
rect 12633 13685 12667 13719
rect 12817 13685 12851 13719
rect 15669 13685 15703 13719
rect 16773 13685 16807 13719
rect 22385 13685 22419 13719
rect 22826 13685 22860 13719
rect 26433 13685 26467 13719
rect 27629 13685 27663 13719
rect 3801 13481 3835 13515
rect 11621 13481 11655 13515
rect 12081 13481 12115 13515
rect 20453 13481 20487 13515
rect 23489 13481 23523 13515
rect 26341 13481 26375 13515
rect 27537 13481 27571 13515
rect 12541 13413 12575 13447
rect 2605 13345 2639 13379
rect 4445 13345 4479 13379
rect 15025 13345 15059 13379
rect 15301 13345 15335 13379
rect 17049 13345 17083 13379
rect 26157 13345 26191 13379
rect 27905 13345 27939 13379
rect 2053 13277 2087 13311
rect 2697 13277 2731 13311
rect 4261 13277 4295 13311
rect 7665 13277 7699 13311
rect 7941 13277 7975 13311
rect 8217 13277 8251 13311
rect 10517 13277 10551 13311
rect 10609 13277 10643 13311
rect 10793 13277 10827 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11805 13277 11839 13311
rect 11897 13277 11931 13311
rect 12173 13277 12207 13311
rect 12266 13277 12300 13311
rect 13277 13277 13311 13311
rect 13461 13277 13495 13311
rect 17693 13277 17727 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 23397 13277 23431 13311
rect 24133 13277 24167 13311
rect 26433 13277 26467 13311
rect 26985 13277 27019 13311
rect 27261 13277 27295 13311
rect 27629 13277 27663 13311
rect 4169 13209 4203 13243
rect 6285 13209 6319 13243
rect 6469 13209 6503 13243
rect 11621 13209 11655 13243
rect 20913 13209 20947 13243
rect 24409 13209 24443 13243
rect 2145 13141 2179 13175
rect 3065 13141 3099 13175
rect 6101 13141 6135 13175
rect 7481 13141 7515 13175
rect 7849 13141 7883 13175
rect 8125 13141 8159 13175
rect 13645 13141 13679 13175
rect 17785 13141 17819 13175
rect 22385 13141 22419 13175
rect 27169 13141 27203 13175
rect 27353 13141 27387 13175
rect 29377 13141 29411 13175
rect 3525 12937 3559 12971
rect 6009 12937 6043 12971
rect 6745 12937 6779 12971
rect 8309 12937 8343 12971
rect 9045 12937 9079 12971
rect 9873 12937 9907 12971
rect 18429 12937 18463 12971
rect 20913 12937 20947 12971
rect 21925 12937 21959 12971
rect 25053 12937 25087 12971
rect 27537 12937 27571 12971
rect 28825 12937 28859 12971
rect 6653 12869 6687 12903
rect 9321 12869 9355 12903
rect 9413 12869 9447 12903
rect 10057 12869 10091 12903
rect 14841 12869 14875 12903
rect 20545 12869 20579 12903
rect 21281 12869 21315 12903
rect 21373 12869 21407 12903
rect 27629 12869 27663 12903
rect 1409 12801 1443 12835
rect 3893 12801 3927 12835
rect 4261 12801 4295 12835
rect 6561 12801 6595 12835
rect 7205 12801 7239 12835
rect 7389 12801 7423 12835
rect 7481 12801 7515 12835
rect 7573 12801 7607 12835
rect 7757 12801 7791 12835
rect 7849 12801 7883 12835
rect 8217 12801 8251 12835
rect 8493 12801 8527 12835
rect 8769 12801 8803 12835
rect 8861 12801 8895 12835
rect 9137 12801 9171 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10149 12801 10183 12835
rect 10333 12801 10367 12835
rect 11253 12801 11287 12835
rect 14565 12801 14599 12835
rect 16681 12801 16715 12835
rect 18613 12801 18647 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 25421 12801 25455 12835
rect 25881 12801 25915 12835
rect 26617 12801 26651 12835
rect 26801 12801 26835 12835
rect 27077 12801 27111 12835
rect 27169 12801 27203 12835
rect 27261 12801 27295 12835
rect 27813 12801 27847 12835
rect 27997 12801 28031 12835
rect 28917 12801 28951 12835
rect 29285 12801 29319 12835
rect 1685 12733 1719 12767
rect 3433 12733 3467 12767
rect 3985 12733 4019 12767
rect 4537 12733 4571 12767
rect 6929 12733 6963 12767
rect 8585 12733 8619 12767
rect 16957 12733 16991 12767
rect 18889 12733 18923 12767
rect 21557 12733 21591 12767
rect 25513 12733 25547 12767
rect 26065 12733 26099 12767
rect 26709 12733 26743 12767
rect 27353 12733 27387 12767
rect 9689 12665 9723 12699
rect 29101 12665 29135 12699
rect 6377 12597 6411 12631
rect 7389 12597 7423 12631
rect 8033 12597 8067 12631
rect 10057 12597 10091 12631
rect 10149 12597 10183 12631
rect 11161 12597 11195 12631
rect 16313 12597 16347 12631
rect 20361 12597 20395 12631
rect 25697 12597 25731 12631
rect 1869 12393 1903 12427
rect 5273 12393 5307 12427
rect 6009 12393 6043 12427
rect 6193 12393 6227 12427
rect 6561 12393 6595 12427
rect 7665 12393 7699 12427
rect 9597 12393 9631 12427
rect 10057 12393 10091 12427
rect 10517 12393 10551 12427
rect 11345 12393 11379 12427
rect 11529 12393 11563 12427
rect 12633 12393 12667 12427
rect 14473 12393 14507 12427
rect 14657 12393 14691 12427
rect 15761 12393 15795 12427
rect 17233 12393 17267 12427
rect 19257 12393 19291 12427
rect 27169 12393 27203 12427
rect 10241 12325 10275 12359
rect 14105 12325 14139 12359
rect 15117 12325 15151 12359
rect 2513 12257 2547 12291
rect 3801 12257 3835 12291
rect 4077 12257 4111 12291
rect 7849 12257 7883 12291
rect 17785 12257 17819 12291
rect 19901 12257 19935 12291
rect 22385 12257 22419 12291
rect 23121 12257 23155 12291
rect 24961 12257 24995 12291
rect 25697 12257 25731 12291
rect 1501 12189 1535 12223
rect 2329 12189 2363 12223
rect 4169 12189 4203 12223
rect 5181 12189 5215 12223
rect 6469 12189 6503 12223
rect 6653 12189 6687 12223
rect 7573 12189 7607 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 9781 12189 9815 12223
rect 9873 12189 9907 12223
rect 10149 12189 10183 12223
rect 10425 12189 10459 12223
rect 10517 12189 10551 12223
rect 10793 12189 10827 12223
rect 11069 12189 11103 12223
rect 11161 12189 11195 12223
rect 11437 12189 11471 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 13093 12189 13127 12223
rect 13277 12189 13311 12223
rect 14933 12189 14967 12223
rect 15853 12189 15887 12223
rect 19717 12189 19751 12223
rect 21833 12189 21867 12223
rect 22017 12189 22051 12223
rect 22293 12189 22327 12223
rect 22477 12189 22511 12223
rect 23213 12189 23247 12223
rect 25421 12189 25455 12223
rect 27445 12189 27479 12223
rect 6147 12155 6181 12189
rect 1685 12121 1719 12155
rect 6377 12121 6411 12155
rect 10701 12121 10735 12155
rect 10977 12121 11011 12155
rect 14749 12121 14783 12155
rect 21925 12121 21959 12155
rect 24777 12121 24811 12155
rect 27353 12121 27387 12155
rect 2237 12053 2271 12087
rect 8125 12053 8159 12087
rect 8309 12053 8343 12087
rect 14473 12053 14507 12087
rect 17601 12053 17635 12087
rect 17693 12053 17727 12087
rect 19625 12053 19659 12087
rect 23581 12053 23615 12087
rect 24409 12053 24443 12087
rect 24869 12053 24903 12087
rect 5549 11849 5583 11883
rect 9597 11849 9631 11883
rect 11529 11849 11563 11883
rect 17509 11849 17543 11883
rect 5273 11781 5307 11815
rect 7874 11781 7908 11815
rect 12449 11781 12483 11815
rect 14013 11781 14047 11815
rect 14565 11781 14599 11815
rect 21833 11781 21867 11815
rect 25697 11781 25731 11815
rect 27445 11781 27479 11815
rect 27905 11781 27939 11815
rect 4997 11713 5031 11747
rect 5181 11713 5215 11747
rect 5365 11713 5399 11747
rect 7389 11713 7423 11747
rect 8125 11713 8159 11747
rect 9045 11713 9079 11747
rect 9229 11713 9263 11747
rect 9321 11713 9355 11747
rect 9413 11713 9447 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 10885 11713 10919 11747
rect 11708 11713 11742 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12080 11713 12114 11747
rect 12173 11713 12207 11747
rect 12909 11713 12943 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 13461 11713 13495 11747
rect 13737 11713 13771 11747
rect 13921 11713 13955 11747
rect 14105 11713 14139 11747
rect 14197 11713 14231 11747
rect 14841 11713 14875 11747
rect 15025 11713 15059 11747
rect 17141 11713 17175 11747
rect 19073 11713 19107 11747
rect 19257 11713 19291 11747
rect 20453 11713 20487 11747
rect 21005 11713 21039 11747
rect 23397 11713 23431 11747
rect 23673 11713 23707 11747
rect 25789 11713 25823 11747
rect 27353 11713 27387 11747
rect 27537 11713 27571 11747
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 12817 11645 12851 11679
rect 13645 11645 13679 11679
rect 17233 11645 17267 11679
rect 20545 11645 20579 11679
rect 20821 11645 20855 11679
rect 23949 11645 23983 11679
rect 27629 11645 27663 11679
rect 8033 11577 8067 11611
rect 11069 11577 11103 11611
rect 13093 11577 13127 11611
rect 14933 11577 14967 11611
rect 8217 11509 8251 11543
rect 12541 11509 12575 11543
rect 14565 11509 14599 11543
rect 14749 11509 14783 11543
rect 19257 11509 19291 11543
rect 25421 11509 25455 11543
rect 29377 11509 29411 11543
rect 1869 11305 1903 11339
rect 2513 11305 2547 11339
rect 4445 11305 4479 11339
rect 6193 11305 6227 11339
rect 9689 11305 9723 11339
rect 10609 11305 10643 11339
rect 11621 11305 11655 11339
rect 14914 11305 14948 11339
rect 16405 11305 16439 11339
rect 19717 11305 19751 11339
rect 21557 11305 21591 11339
rect 22845 11305 22879 11339
rect 23029 11305 23063 11339
rect 28089 11305 28123 11339
rect 28825 11305 28859 11339
rect 10517 11237 10551 11271
rect 19625 11237 19659 11271
rect 19809 11237 19843 11271
rect 21281 11237 21315 11271
rect 27997 11237 28031 11271
rect 29193 11237 29227 11271
rect 1685 11169 1719 11203
rect 2329 11169 2363 11203
rect 3801 11169 3835 11203
rect 4077 11169 4111 11203
rect 4537 11169 4571 11203
rect 4813 11169 4847 11203
rect 6285 11169 6319 11203
rect 10701 11169 10735 11203
rect 11713 11169 11747 11203
rect 11805 11169 11839 11203
rect 18797 11169 18831 11203
rect 22017 11169 22051 11203
rect 22293 11169 22327 11203
rect 22753 11169 22787 11203
rect 23213 11169 23247 11203
rect 1593 11101 1627 11135
rect 2237 11101 2271 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2789 11101 2823 11135
rect 3157 11101 3191 11135
rect 4169 11101 4203 11135
rect 4905 11101 4939 11135
rect 6193 11101 6227 11135
rect 6469 11101 6503 11135
rect 7021 11101 7055 11135
rect 9137 11101 9171 11135
rect 9321 11101 9355 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 10425 11101 10459 11135
rect 11897 11101 11931 11135
rect 12081 11101 12115 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 13001 11101 13035 11135
rect 13093 11101 13127 11135
rect 14657 11101 14691 11135
rect 16681 11101 16715 11135
rect 17049 11101 17083 11135
rect 17233 11101 17267 11135
rect 17325 11101 17359 11135
rect 17509 11101 17543 11135
rect 17601 11101 17635 11135
rect 17785 11101 17819 11135
rect 18705 11101 18739 11135
rect 18889 11101 18923 11135
rect 19993 11101 20027 11135
rect 20269 11101 20303 11135
rect 20545 11101 20579 11135
rect 20637 11101 20671 11135
rect 20821 11101 20855 11135
rect 20913 11101 20947 11135
rect 21005 11101 21039 11135
rect 21373 11101 21407 11135
rect 21557 11101 21591 11135
rect 22109 11101 22143 11135
rect 22385 11101 22419 11135
rect 23029 11101 23063 11135
rect 23305 11101 23339 11135
rect 26065 11101 26099 11135
rect 26341 11101 26375 11135
rect 27629 11101 27663 11135
rect 28089 11101 28123 11135
rect 28273 11101 28307 11135
rect 28917 11101 28951 11135
rect 29377 11101 29411 11135
rect 2881 11033 2915 11067
rect 3019 11033 3053 11067
rect 3433 11033 3467 11067
rect 3617 11033 3651 11067
rect 4286 11033 4320 11067
rect 9229 11033 9263 11067
rect 11529 11033 11563 11067
rect 16589 11033 16623 11067
rect 17693 11033 17727 11067
rect 19257 11033 19291 11067
rect 20361 11033 20395 11067
rect 21281 11033 21315 11067
rect 21649 11033 21683 11067
rect 21833 11033 21867 11067
rect 26249 11033 26283 11067
rect 27445 11033 27479 11067
rect 27721 11033 27755 11067
rect 3249 10965 3283 10999
rect 6653 10965 6687 10999
rect 8309 10965 8343 10999
rect 8953 10965 8987 10999
rect 12909 10965 12943 10999
rect 13185 10965 13219 10999
rect 17141 10965 17175 10999
rect 17417 10965 17451 10999
rect 20177 10965 20211 10999
rect 21097 10965 21131 10999
rect 25973 10965 26007 10999
rect 27813 10965 27847 10999
rect 3525 10761 3559 10795
rect 7113 10761 7147 10795
rect 8125 10761 8159 10795
rect 14105 10761 14139 10795
rect 18889 10761 18923 10795
rect 19165 10761 19199 10795
rect 19701 10761 19735 10795
rect 20085 10761 20119 10795
rect 21097 10761 21131 10795
rect 21925 10761 21959 10795
rect 26801 10761 26835 10795
rect 1501 10693 1535 10727
rect 3617 10693 3651 10727
rect 6745 10693 6779 10727
rect 10609 10693 10643 10727
rect 13277 10693 13311 10727
rect 13369 10693 13403 10727
rect 13921 10693 13955 10727
rect 17969 10693 18003 10727
rect 19901 10693 19935 10727
rect 20453 10693 20487 10727
rect 25329 10693 25363 10727
rect 27537 10693 27571 10727
rect 27753 10693 27787 10727
rect 1685 10625 1719 10659
rect 2605 10625 2639 10659
rect 2789 10625 2823 10659
rect 2973 10625 3007 10659
rect 3065 10625 3099 10659
rect 3801 10625 3835 10659
rect 3985 10625 4019 10659
rect 5089 10625 5123 10659
rect 5457 10625 5491 10659
rect 6929 10625 6963 10659
rect 7389 10625 7423 10659
rect 8401 10625 8435 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 9413 10625 9447 10659
rect 9597 10625 9631 10659
rect 10425 10625 10459 10659
rect 10701 10625 10735 10659
rect 10793 10625 10827 10659
rect 13553 10625 13587 10659
rect 13645 10625 13679 10659
rect 13737 10625 13771 10659
rect 14013 10625 14047 10659
rect 16773 10625 16807 10659
rect 16957 10625 16991 10659
rect 17233 10625 17267 10659
rect 17417 10625 17451 10659
rect 17877 10625 17911 10659
rect 18797 10625 18831 10659
rect 18981 10625 19015 10659
rect 19073 10625 19107 10659
rect 19257 10625 19291 10659
rect 20269 10625 20303 10659
rect 21281 10625 21315 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22845 10625 22879 10659
rect 27997 10625 28031 10659
rect 28181 10625 28215 10659
rect 5365 10557 5399 10591
rect 5733 10557 5767 10591
rect 16865 10557 16899 10591
rect 21465 10557 21499 10591
rect 23121 10557 23155 10591
rect 24869 10557 24903 10591
rect 25053 10557 25087 10591
rect 3341 10489 3375 10523
rect 5273 10489 5307 10523
rect 5549 10489 5583 10523
rect 19533 10489 19567 10523
rect 27905 10489 27939 10523
rect 4905 10421 4939 10455
rect 5457 10421 5491 10455
rect 8309 10421 8343 10455
rect 8769 10421 8803 10455
rect 9413 10421 9447 10455
rect 10977 10421 11011 10455
rect 11805 10421 11839 10455
rect 17417 10421 17451 10455
rect 19717 10421 19751 10455
rect 27721 10421 27755 10455
rect 27997 10421 28031 10455
rect 4169 10217 4203 10251
rect 6377 10217 6411 10251
rect 7021 10217 7055 10251
rect 7665 10217 7699 10251
rect 7941 10217 7975 10251
rect 9689 10217 9723 10251
rect 10793 10217 10827 10251
rect 12817 10217 12851 10251
rect 13737 10217 13771 10251
rect 13921 10217 13955 10251
rect 15681 10217 15715 10251
rect 16589 10217 16623 10251
rect 17509 10217 17543 10251
rect 18153 10217 18187 10251
rect 19533 10217 19567 10251
rect 19717 10217 19751 10251
rect 20085 10217 20119 10251
rect 22845 10217 22879 10251
rect 24133 10217 24167 10251
rect 27537 10217 27571 10251
rect 6837 10149 6871 10183
rect 12725 10149 12759 10183
rect 14197 10149 14231 10183
rect 17693 10149 17727 10183
rect 6745 10081 6779 10115
rect 15945 10081 15979 10115
rect 16313 10081 16347 10115
rect 19349 10081 19383 10115
rect 21649 10081 21683 10115
rect 23305 10081 23339 10115
rect 23489 10081 23523 10115
rect 26065 10081 26099 10115
rect 26341 10081 26375 10115
rect 27629 10081 27663 10115
rect 27905 10081 27939 10115
rect 4353 10013 4387 10047
rect 4629 10013 4663 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 6561 10013 6595 10047
rect 7849 10013 7883 10047
rect 8033 10013 8067 10047
rect 9873 10013 9907 10047
rect 9965 10013 9999 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 10609 10013 10643 10047
rect 10885 10013 10919 10047
rect 11805 10013 11839 10047
rect 12817 10013 12851 10047
rect 13277 10013 13311 10047
rect 16221 10013 16255 10047
rect 18337 10013 18371 10047
rect 18521 10013 18555 10047
rect 18705 10013 18739 10047
rect 19533 10013 19567 10047
rect 19993 10013 20027 10047
rect 21741 10013 21775 10047
rect 24225 10013 24259 10047
rect 25973 10013 26007 10047
rect 27261 10013 27295 10047
rect 7205 9945 7239 9979
rect 12541 9945 12575 9979
rect 13093 9945 13127 9979
rect 13553 9945 13587 9979
rect 17325 9945 17359 9979
rect 18429 9945 18463 9979
rect 19257 9945 19291 9979
rect 23213 9945 23247 9979
rect 27353 9945 27387 9979
rect 27537 9945 27571 9979
rect 4537 9877 4571 9911
rect 4997 9877 5031 9911
rect 7005 9877 7039 9911
rect 10333 9877 10367 9911
rect 13461 9877 13495 9911
rect 13753 9877 13787 9911
rect 17535 9877 17569 9911
rect 22109 9877 22143 9911
rect 29377 9877 29411 9911
rect 4905 9673 4939 9707
rect 8861 9673 8895 9707
rect 10149 9673 10183 9707
rect 13737 9673 13771 9707
rect 21373 9673 21407 9707
rect 4997 9605 5031 9639
rect 9387 9605 9421 9639
rect 11989 9605 12023 9639
rect 14933 9605 14967 9639
rect 21925 9605 21959 9639
rect 23673 9605 23707 9639
rect 27261 9605 27295 9639
rect 29009 9605 29043 9639
rect 3893 9537 3927 9571
rect 6929 9537 6963 9571
rect 7113 9537 7147 9571
rect 7389 9537 7423 9571
rect 7481 9537 7515 9571
rect 8777 9537 8811 9571
rect 9262 9537 9296 9571
rect 9781 9537 9815 9571
rect 9873 9537 9907 9571
rect 9965 9537 9999 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 13645 9537 13679 9571
rect 13829 9537 13863 9571
rect 15025 9537 15059 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 17509 9537 17543 9571
rect 20913 9537 20947 9571
rect 21097 9537 21131 9571
rect 21281 9537 21315 9571
rect 21465 9537 21499 9571
rect 21833 9537 21867 9571
rect 22017 9537 22051 9571
rect 23489 9537 23523 9571
rect 23581 9537 23615 9571
rect 23857 9537 23891 9571
rect 29101 9537 29135 9571
rect 29193 9537 29227 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 5181 9469 5215 9503
rect 9689 9469 9723 9503
rect 10149 9469 10183 9503
rect 11621 9469 11655 9503
rect 16957 9469 16991 9503
rect 21005 9469 21039 9503
rect 26985 9469 27019 9503
rect 28733 9469 28767 9503
rect 7205 9401 7239 9435
rect 29377 9401 29411 9435
rect 3525 9333 3559 9367
rect 4537 9333 4571 9367
rect 6653 9333 6687 9367
rect 6929 9333 6963 9367
rect 9137 9333 9171 9367
rect 12173 9333 12207 9367
rect 16773 9333 16807 9367
rect 17509 9333 17543 9367
rect 23305 9333 23339 9367
rect 2145 9129 2179 9163
rect 2329 9129 2363 9163
rect 6653 9129 6687 9163
rect 8677 9129 8711 9163
rect 10609 9129 10643 9163
rect 13369 9129 13403 9163
rect 16957 9129 16991 9163
rect 23029 9129 23063 9163
rect 27353 9129 27387 9163
rect 9413 9061 9447 9095
rect 19257 9061 19291 9095
rect 22385 9061 22419 9095
rect 2789 8993 2823 9027
rect 2973 8993 3007 9027
rect 4261 8993 4295 9027
rect 6377 8993 6411 9027
rect 9873 8993 9907 9027
rect 10057 8993 10091 9027
rect 12173 8993 12207 9027
rect 13277 8993 13311 9027
rect 13645 8993 13679 9027
rect 13737 8993 13771 9027
rect 15853 8993 15887 9027
rect 17785 8993 17819 9027
rect 21005 8993 21039 9027
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 3985 8925 4019 8959
rect 6285 8925 6319 8959
rect 6929 8925 6963 8959
rect 9137 8925 9171 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 10333 8925 10367 8959
rect 10425 8925 10459 8959
rect 10517 8925 10551 8959
rect 10793 8925 10827 8959
rect 11069 8925 11103 8959
rect 11162 8925 11196 8959
rect 11437 8925 11471 8959
rect 11575 8925 11609 8959
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 12817 8925 12851 8959
rect 12909 8925 12943 8959
rect 13001 8925 13035 8959
rect 13553 8925 13587 8959
rect 13829 8925 13863 8959
rect 15577 8925 15611 8959
rect 17141 8925 17175 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 17877 8925 17911 8959
rect 21097 8925 21131 8959
rect 22109 8925 22143 8959
rect 22661 8925 22695 8959
rect 23208 8925 23242 8959
rect 23397 8925 23431 8959
rect 23525 8925 23559 8959
rect 23673 8925 23707 8959
rect 24501 8925 24535 8959
rect 27261 8925 27295 8959
rect 6009 8857 6043 8891
rect 7205 8857 7239 8891
rect 9045 8857 9079 8891
rect 10701 8857 10735 8891
rect 10885 8857 10919 8891
rect 11345 8857 11379 8891
rect 12541 8857 12575 8891
rect 20729 8857 20763 8891
rect 22753 8857 22787 8891
rect 23305 8857 23339 8891
rect 10241 8789 10275 8823
rect 11713 8789 11747 8823
rect 15209 8789 15243 8823
rect 15669 8789 15703 8823
rect 18245 8789 18279 8823
rect 21189 8789 21223 8823
rect 22569 8789 22603 8823
rect 24593 8789 24627 8823
rect 5089 8585 5123 8619
rect 6929 8585 6963 8619
rect 11621 8585 11655 8619
rect 12639 8585 12673 8619
rect 13921 8585 13955 8619
rect 16221 8585 16255 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 19257 8585 19291 8619
rect 19625 8585 19659 8619
rect 20085 8585 20119 8619
rect 23397 8585 23431 8619
rect 24133 8585 24167 8619
rect 29193 8585 29227 8619
rect 7573 8517 7607 8551
rect 12541 8517 12575 8551
rect 14749 8517 14783 8551
rect 16405 8517 16439 8551
rect 1685 8449 1719 8483
rect 4997 8449 5031 8483
rect 7205 8449 7239 8483
rect 11713 8449 11747 8483
rect 12725 8449 12759 8483
rect 12817 8449 12851 8483
rect 13829 8449 13863 8483
rect 14013 8449 14047 8483
rect 14473 8449 14507 8483
rect 16497 8449 16531 8483
rect 16957 8449 16991 8483
rect 17141 8449 17175 8483
rect 17325 8449 17359 8483
rect 17509 8449 17543 8483
rect 19165 8449 19199 8483
rect 20177 8449 20211 8483
rect 20269 8449 20303 8483
rect 20362 8449 20396 8483
rect 23581 8449 23615 8483
rect 23673 8449 23707 8483
rect 23949 8449 23983 8483
rect 24041 8449 24075 8483
rect 25697 8449 25731 8483
rect 29285 8449 29319 8483
rect 1409 8381 1443 8415
rect 7113 8381 7147 8415
rect 7481 8381 7515 8415
rect 18981 8381 19015 8415
rect 23857 8313 23891 8347
rect 25605 8313 25639 8347
rect 20453 8245 20487 8279
rect 6285 8041 6319 8075
rect 10333 8041 10367 8075
rect 11437 8041 11471 8075
rect 12265 8041 12299 8075
rect 13829 8041 13863 8075
rect 15577 8041 15611 8075
rect 4721 7973 4755 8007
rect 10977 7973 11011 8007
rect 21833 7973 21867 8007
rect 22017 7973 22051 8007
rect 1685 7905 1719 7939
rect 3065 7905 3099 7939
rect 3341 7905 3375 7939
rect 4997 7905 5031 7939
rect 5917 7905 5951 7939
rect 6009 7905 6043 7939
rect 9689 7905 9723 7939
rect 21005 7905 21039 7939
rect 23765 7905 23799 7939
rect 1409 7837 1443 7871
rect 2973 7837 3007 7871
rect 5089 7837 5123 7871
rect 5641 7837 5675 7871
rect 6837 7837 6871 7871
rect 7113 7837 7147 7871
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 10517 7837 10551 7871
rect 10609 7837 10643 7871
rect 10885 7837 10919 7871
rect 11161 7837 11195 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 13001 7837 13035 7871
rect 13093 7837 13127 7871
rect 13461 7837 13495 7871
rect 13645 7837 13679 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14289 7837 14323 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 14657 7837 14691 7871
rect 15485 7837 15519 7871
rect 17233 7837 17267 7871
rect 19533 7837 19567 7871
rect 19717 7837 19751 7871
rect 19809 7837 19843 7871
rect 20361 7837 20395 7871
rect 20453 7837 20487 7871
rect 20545 7837 20579 7871
rect 20729 7837 20763 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21281 7837 21315 7871
rect 22288 7837 22322 7871
rect 22385 7837 22419 7871
rect 22660 7837 22694 7871
rect 22753 7837 22787 7871
rect 23121 7837 23155 7871
rect 23397 7837 23431 7871
rect 23489 7837 23523 7871
rect 23949 7837 23983 7871
rect 24225 7837 24259 7871
rect 24593 7837 24627 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 29377 7837 29411 7871
rect 6126 7769 6160 7803
rect 7021 7769 7055 7803
rect 10701 7769 10735 7803
rect 12081 7769 12115 7803
rect 14841 7769 14875 7803
rect 21465 7769 21499 7803
rect 21557 7769 21591 7803
rect 22477 7769 22511 7803
rect 23305 7769 23339 7803
rect 24777 7769 24811 7803
rect 6653 7701 6687 7735
rect 8033 7701 8067 7735
rect 8309 7701 8343 7735
rect 13553 7701 13587 7735
rect 17141 7701 17175 7735
rect 19349 7701 19383 7735
rect 20177 7701 20211 7735
rect 22109 7701 22143 7735
rect 23673 7701 23707 7735
rect 24133 7701 24167 7735
rect 24409 7701 24443 7735
rect 29193 7701 29227 7735
rect 2881 7497 2915 7531
rect 3341 7497 3375 7531
rect 6653 7497 6687 7531
rect 12265 7497 12299 7531
rect 12357 7497 12391 7531
rect 14473 7497 14507 7531
rect 15945 7497 15979 7531
rect 16865 7497 16899 7531
rect 20085 7497 20119 7531
rect 22385 7497 22419 7531
rect 22477 7497 22511 7531
rect 24593 7497 24627 7531
rect 4077 7429 4111 7463
rect 5457 7429 5491 7463
rect 7205 7429 7239 7463
rect 7573 7429 7607 7463
rect 9597 7429 9631 7463
rect 14197 7429 14231 7463
rect 18429 7429 18463 7463
rect 21189 7429 21223 7463
rect 21281 7429 21315 7463
rect 3709 7361 3743 7395
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 4905 7361 4939 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 5979 7361 6013 7395
rect 6837 7361 6871 7395
rect 7113 7361 7147 7395
rect 7389 7361 7423 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 8309 7361 8343 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 9229 7361 9263 7395
rect 9689 7361 9723 7395
rect 9781 7361 9815 7395
rect 10149 7361 10183 7395
rect 10609 7361 10643 7395
rect 10977 7361 11011 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 11897 7361 11931 7395
rect 12081 7361 12115 7395
rect 12541 7361 12575 7395
rect 12909 7361 12943 7395
rect 13093 7361 13127 7395
rect 13829 7361 13863 7395
rect 13922 7361 13956 7395
rect 14105 7361 14139 7395
rect 14335 7361 14369 7395
rect 15669 7361 15703 7395
rect 16806 7361 16840 7395
rect 17601 7361 17635 7395
rect 17693 7361 17727 7395
rect 17785 7361 17819 7395
rect 17969 7361 18003 7395
rect 19349 7361 19383 7395
rect 19441 7361 19475 7395
rect 19717 7361 19751 7395
rect 20269 7361 20303 7395
rect 20361 7361 20395 7395
rect 20637 7361 20671 7395
rect 21097 7361 21131 7395
rect 21465 7361 21499 7395
rect 22017 7361 22051 7395
rect 22110 7361 22144 7395
rect 22752 7361 22786 7395
rect 22845 7361 22879 7395
rect 24041 7361 24075 7395
rect 24317 7361 24351 7395
rect 24409 7361 24443 7395
rect 2973 7293 3007 7327
rect 3157 7293 3191 7327
rect 3801 7293 3835 7327
rect 4537 7293 4571 7327
rect 5457 7293 5491 7327
rect 5641 7293 5675 7327
rect 7021 7293 7055 7327
rect 9045 7293 9079 7327
rect 9413 7293 9447 7327
rect 10701 7293 10735 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 15301 7293 15335 7327
rect 15761 7293 15795 7327
rect 17325 7293 17359 7327
rect 18613 7293 18647 7327
rect 18705 7293 18739 7327
rect 19073 7293 19107 7327
rect 19165 7293 19199 7327
rect 24133 7293 24167 7327
rect 4445 7225 4479 7259
rect 6193 7225 6227 7259
rect 8861 7225 8895 7259
rect 10517 7225 10551 7259
rect 16681 7225 16715 7259
rect 20913 7225 20947 7259
rect 2513 7157 2547 7191
rect 4629 7157 4663 7191
rect 7113 7157 7147 7191
rect 7757 7157 7791 7191
rect 8401 7157 8435 7191
rect 9873 7157 9907 7191
rect 17233 7157 17267 7191
rect 17417 7157 17451 7191
rect 19625 7157 19659 7191
rect 20545 7157 20579 7191
rect 1672 6953 1706 6987
rect 3157 6953 3191 6987
rect 8217 6953 8251 6987
rect 8953 6953 8987 6987
rect 10149 6953 10183 6987
rect 12725 6953 12759 6987
rect 15301 6953 15335 6987
rect 18889 6953 18923 6987
rect 12633 6885 12667 6919
rect 1409 6817 1443 6851
rect 4537 6817 4571 6851
rect 7849 6817 7883 6851
rect 10609 6817 10643 6851
rect 13001 6817 13035 6851
rect 13093 6817 13127 6851
rect 13461 6817 13495 6851
rect 15761 6817 15795 6851
rect 16313 6817 16347 6851
rect 18521 6817 18555 6851
rect 4445 6749 4479 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 12081 6749 12115 6783
rect 12449 6749 12483 6783
rect 12909 6749 12943 6783
rect 13185 6749 13219 6783
rect 13369 6749 13403 6783
rect 13645 6749 13679 6783
rect 13829 6749 13863 6783
rect 15485 6749 15519 6783
rect 15577 6749 15611 6783
rect 15853 6749 15887 6783
rect 16221 6749 16255 6783
rect 16957 6749 16991 6783
rect 17509 6749 17543 6783
rect 17785 6749 17819 6783
rect 18061 6749 18095 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 18797 6749 18831 6783
rect 18981 6749 19015 6783
rect 19441 6749 19475 6783
rect 19809 6749 19843 6783
rect 21189 6749 21223 6783
rect 12265 6681 12299 6715
rect 12357 6681 12391 6715
rect 16773 6681 16807 6715
rect 17693 6681 17727 6715
rect 19533 6681 19567 6715
rect 19625 6681 19659 6715
rect 4813 6613 4847 6647
rect 13737 6613 13771 6647
rect 17141 6613 17175 6647
rect 17325 6613 17359 6647
rect 19257 6613 19291 6647
rect 21097 6613 21131 6647
rect 2421 6409 2455 6443
rect 8125 6409 8159 6443
rect 12633 6409 12667 6443
rect 13369 6409 13403 6443
rect 22385 6409 22419 6443
rect 8401 6341 8435 6375
rect 10241 6341 10275 6375
rect 11805 6341 11839 6375
rect 11897 6341 11931 6375
rect 17141 6341 17175 6375
rect 17233 6341 17267 6375
rect 20361 6341 20395 6375
rect 21189 6341 21223 6375
rect 21281 6341 21315 6375
rect 24041 6341 24075 6375
rect 1409 6273 1443 6307
rect 2329 6273 2363 6307
rect 6561 6273 6595 6307
rect 8309 6273 8343 6307
rect 8493 6273 8527 6307
rect 8677 6273 8711 6307
rect 9965 6273 9999 6307
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 11713 6273 11747 6307
rect 12081 6273 12115 6307
rect 12449 6273 12483 6307
rect 13553 6273 13587 6307
rect 13737 6273 13771 6307
rect 13921 6273 13955 6307
rect 14105 6273 14139 6307
rect 14657 6273 14691 6307
rect 14749 6273 14783 6307
rect 15025 6273 15059 6307
rect 15301 6273 15335 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 17049 6273 17083 6307
rect 17417 6273 17451 6307
rect 20131 6273 20165 6307
rect 20269 6273 20303 6307
rect 20499 6273 20533 6307
rect 20637 6273 20671 6307
rect 21092 6273 21126 6307
rect 21464 6273 21498 6307
rect 21557 6273 21591 6307
rect 21833 6273 21867 6307
rect 22109 6273 22143 6307
rect 22201 6273 22235 6307
rect 22661 6273 22695 6307
rect 22845 6273 22879 6307
rect 22937 6273 22971 6307
rect 23029 6273 23063 6307
rect 23305 6271 23339 6305
rect 23489 6273 23523 6307
rect 23673 6273 23707 6307
rect 23857 6273 23891 6307
rect 24133 6273 24167 6307
rect 24317 6273 24351 6307
rect 24409 6273 24443 6307
rect 24501 6273 24535 6307
rect 24777 6273 24811 6307
rect 25053 6273 25087 6307
rect 25145 6273 25179 6307
rect 29101 6273 29135 6307
rect 1685 6205 1719 6239
rect 6653 6205 6687 6239
rect 12265 6205 12299 6239
rect 13829 6205 13863 6239
rect 15485 6205 15519 6239
rect 15577 6205 15611 6239
rect 23581 6205 23615 6239
rect 29377 6205 29411 6239
rect 6929 6137 6963 6171
rect 15117 6137 15151 6171
rect 21925 6137 21959 6171
rect 23213 6137 23247 6171
rect 24869 6137 24903 6171
rect 10517 6069 10551 6103
rect 11529 6069 11563 6103
rect 14473 6069 14507 6103
rect 14933 6069 14967 6103
rect 16865 6069 16899 6103
rect 19993 6069 20027 6103
rect 20913 6069 20947 6103
rect 24685 6069 24719 6103
rect 25329 6069 25363 6103
rect 8309 5865 8343 5899
rect 11161 5865 11195 5899
rect 11529 5865 11563 5899
rect 13553 5865 13587 5899
rect 16129 5865 16163 5899
rect 18889 5865 18923 5899
rect 19809 5865 19843 5899
rect 22569 5865 22603 5899
rect 8125 5797 8159 5831
rect 8677 5797 8711 5831
rect 8953 5797 8987 5831
rect 10609 5797 10643 5831
rect 14197 5797 14231 5831
rect 21097 5797 21131 5831
rect 7205 5729 7239 5763
rect 8769 5729 8803 5763
rect 16497 5729 16531 5763
rect 16589 5729 16623 5763
rect 17877 5729 17911 5763
rect 21649 5729 21683 5763
rect 4169 5661 4203 5695
rect 7021 5661 7055 5695
rect 7113 5661 7147 5695
rect 8033 5661 8067 5695
rect 8493 5661 8527 5695
rect 9137 5661 9171 5695
rect 9229 5661 9263 5695
rect 9505 5661 9539 5695
rect 10057 5661 10091 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 10885 5661 10919 5695
rect 10977 5661 11011 5695
rect 11253 5661 11287 5695
rect 11713 5661 11747 5695
rect 11897 5661 11931 5695
rect 11989 5661 12023 5695
rect 12909 5661 12943 5695
rect 13057 5661 13091 5695
rect 13415 5661 13449 5695
rect 14381 5661 14415 5695
rect 14565 5661 14599 5695
rect 14657 5661 14691 5695
rect 16313 5661 16347 5695
rect 16681 5661 16715 5695
rect 16865 5661 16899 5695
rect 17233 5661 17267 5695
rect 17417 5661 17451 5695
rect 17601 5661 17635 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 18337 5661 18371 5695
rect 18429 5661 18463 5695
rect 18613 5661 18647 5695
rect 18705 5661 18739 5695
rect 18981 5661 19015 5695
rect 19717 5661 19751 5695
rect 19993 5661 20027 5695
rect 20085 5661 20119 5695
rect 20637 5661 20671 5695
rect 20913 5661 20947 5695
rect 21097 5661 21131 5695
rect 21189 5661 21223 5695
rect 21373 5661 21407 5695
rect 21741 5661 21775 5695
rect 22753 5661 22787 5695
rect 22937 5661 22971 5695
rect 24593 5661 24627 5695
rect 24777 5661 24811 5695
rect 24961 5661 24995 5695
rect 4445 5593 4479 5627
rect 9321 5593 9355 5627
rect 10241 5593 10275 5627
rect 13185 5593 13219 5627
rect 13277 5593 13311 5627
rect 17509 5593 17543 5627
rect 24685 5593 24719 5627
rect 5917 5525 5951 5559
rect 6653 5525 6687 5559
rect 10701 5525 10735 5559
rect 17785 5525 17819 5559
rect 20269 5525 20303 5559
rect 20729 5525 20763 5559
rect 21373 5525 21407 5559
rect 24409 5525 24443 5559
rect 4721 5321 4755 5355
rect 5089 5321 5123 5355
rect 5641 5321 5675 5355
rect 8125 5321 8159 5355
rect 8769 5321 8803 5355
rect 10057 5321 10091 5355
rect 11529 5321 11563 5355
rect 12725 5321 12759 5355
rect 14105 5321 14139 5355
rect 14933 5321 14967 5355
rect 16497 5321 16531 5355
rect 16865 5321 16899 5355
rect 18153 5321 18187 5355
rect 20453 5321 20487 5355
rect 22109 5321 22143 5355
rect 23949 5321 23983 5355
rect 5181 5253 5215 5287
rect 6653 5253 6687 5287
rect 8309 5253 8343 5287
rect 10425 5253 10459 5287
rect 10885 5253 10919 5287
rect 14197 5253 14231 5287
rect 14565 5253 14599 5287
rect 17785 5253 17819 5287
rect 18613 5253 18647 5287
rect 22385 5253 22419 5287
rect 1501 5185 1535 5219
rect 5733 5185 5767 5219
rect 8401 5185 8435 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 9321 5185 9355 5219
rect 10241 5185 10275 5219
rect 10517 5185 10551 5219
rect 11069 5185 11103 5219
rect 11253 5185 11287 5219
rect 11345 5185 11379 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12081 5185 12115 5219
rect 12909 5185 12943 5219
rect 13001 5185 13035 5219
rect 13093 5185 13127 5219
rect 13277 5185 13311 5219
rect 13369 5185 13403 5219
rect 13553 5185 13587 5219
rect 13921 5185 13955 5219
rect 14381 5185 14415 5219
rect 14657 5185 14691 5219
rect 15117 5185 15151 5219
rect 15209 5185 15243 5219
rect 15485 5185 15519 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 16221 5185 16255 5219
rect 16313 5185 16347 5219
rect 16681 5185 16715 5219
rect 16865 5185 16899 5219
rect 17141 5185 17175 5219
rect 17325 5185 17359 5219
rect 17417 5185 17451 5219
rect 17509 5185 17543 5219
rect 17969 5185 18003 5219
rect 18245 5185 18279 5219
rect 18797 5185 18831 5219
rect 18889 5185 18923 5219
rect 19165 5185 19199 5219
rect 19441 5185 19475 5219
rect 19533 5185 19567 5219
rect 20085 5185 20119 5219
rect 20269 5185 20303 5219
rect 20545 5185 20579 5219
rect 20913 5185 20947 5219
rect 21097 5185 21131 5219
rect 21189 5185 21223 5219
rect 21465 5185 21499 5219
rect 22247 5185 22281 5219
rect 22477 5185 22511 5219
rect 22660 5185 22694 5219
rect 22753 5185 22787 5219
rect 24041 5185 24075 5219
rect 29285 5185 29319 5219
rect 5365 5117 5399 5151
rect 6377 5117 6411 5151
rect 13645 5117 13679 5151
rect 13737 5117 13771 5151
rect 19257 5117 19291 5151
rect 9229 5049 9263 5083
rect 15393 5049 15427 5083
rect 17693 5049 17727 5083
rect 19073 5049 19107 5083
rect 29101 5049 29135 5083
rect 1593 4981 1627 5015
rect 11989 4981 12023 5015
rect 21373 4981 21407 5015
rect 13829 4777 13863 4811
rect 14841 4777 14875 4811
rect 15301 4777 15335 4811
rect 16865 4777 16899 4811
rect 18521 4777 18555 4811
rect 22385 4777 22419 4811
rect 23949 4777 23983 4811
rect 11989 4709 12023 4743
rect 18981 4709 19015 4743
rect 22293 4709 22327 4743
rect 22477 4709 22511 4743
rect 22937 4709 22971 4743
rect 21925 4641 21959 4675
rect 23397 4641 23431 4675
rect 11529 4573 11563 4607
rect 11713 4573 11747 4607
rect 11897 4573 11931 4607
rect 12725 4573 12759 4607
rect 13277 4573 13311 4607
rect 13461 4573 13495 4607
rect 13645 4573 13679 4607
rect 15025 4573 15059 4607
rect 15117 4573 15151 4607
rect 15393 4573 15427 4607
rect 16773 4573 16807 4607
rect 18705 4573 18739 4607
rect 18797 4573 18831 4607
rect 19073 4573 19107 4607
rect 20361 4573 20395 4607
rect 22691 4573 22725 4607
rect 22845 4573 22879 4607
rect 23151 4573 23185 4607
rect 23305 4573 23339 4607
rect 23581 4573 23615 4607
rect 24041 4573 24075 4607
rect 24501 4573 24535 4607
rect 12817 4505 12851 4539
rect 13553 4505 13587 4539
rect 11529 4437 11563 4471
rect 20453 4437 20487 4471
rect 23765 4437 23799 4471
rect 24593 4437 24627 4471
rect 10701 4233 10735 4267
rect 12725 4233 12759 4267
rect 15117 4233 15151 4267
rect 17785 4233 17819 4267
rect 19165 4233 19199 4267
rect 10977 4165 11011 4199
rect 11161 4165 11195 4199
rect 11713 4165 11747 4199
rect 12541 4165 12575 4199
rect 12817 4165 12851 4199
rect 14749 4165 14783 4199
rect 23765 4165 23799 4199
rect 8953 4097 8987 4131
rect 12173 4097 12207 4131
rect 12357 4097 12391 4131
rect 12909 4097 12943 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 15025 4097 15059 4131
rect 16313 4097 16347 4131
rect 16497 4097 16531 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 17693 4097 17727 4131
rect 17969 4097 18003 4131
rect 18153 4097 18187 4131
rect 19073 4097 19107 4131
rect 9229 4029 9263 4063
rect 12265 4029 12299 4063
rect 13277 4029 13311 4063
rect 14381 4029 14415 4063
rect 19441 4029 19475 4063
rect 19717 4029 19751 4063
rect 23489 4029 23523 4063
rect 25237 4029 25271 4063
rect 11345 3961 11379 3995
rect 12081 3961 12115 3995
rect 14933 3961 14967 3995
rect 11529 3893 11563 3927
rect 11713 3893 11747 3927
rect 13093 3893 13127 3927
rect 14749 3893 14783 3927
rect 16405 3893 16439 3927
rect 16681 3893 16715 3927
rect 18061 3893 18095 3927
rect 21189 3893 21223 3927
rect 9965 3689 9999 3723
rect 10701 3689 10735 3723
rect 12725 3689 12759 3723
rect 13461 3689 13495 3723
rect 13645 3689 13679 3723
rect 16589 3689 16623 3723
rect 17969 3689 18003 3723
rect 18705 3689 18739 3723
rect 19809 3689 19843 3723
rect 20269 3689 20303 3723
rect 23121 3689 23155 3723
rect 23305 3689 23339 3723
rect 10333 3621 10367 3655
rect 16221 3621 16255 3655
rect 16773 3621 16807 3655
rect 18429 3621 18463 3655
rect 19993 3621 20027 3655
rect 22477 3621 22511 3655
rect 22569 3621 22603 3655
rect 29101 3621 29135 3655
rect 14381 3553 14415 3587
rect 14657 3553 14691 3587
rect 19441 3553 19475 3587
rect 23857 3553 23891 3587
rect 1501 3485 1535 3519
rect 9873 3485 9907 3519
rect 10977 3485 11011 3519
rect 13001 3485 13035 3519
rect 13185 3485 13219 3519
rect 17693 3485 17727 3519
rect 18245 3485 18279 3519
rect 20453 3485 20487 3519
rect 20729 3485 20763 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 23673 3485 23707 3519
rect 23765 3485 23799 3519
rect 23949 3485 23983 3519
rect 10701 3417 10735 3451
rect 11253 3417 11287 3451
rect 13369 3417 13403 3451
rect 13613 3417 13647 3451
rect 13829 3417 13863 3451
rect 17417 3417 17451 3451
rect 17785 3417 17819 3451
rect 18061 3417 18095 3451
rect 18521 3417 18555 3451
rect 19809 3417 19843 3451
rect 20637 3417 20671 3451
rect 21005 3417 21039 3451
rect 23581 3417 23615 3451
rect 29285 3417 29319 3451
rect 1593 3349 1627 3383
rect 10885 3349 10919 3383
rect 16129 3349 16163 3383
rect 16589 3349 16623 3383
rect 17601 3349 17635 3383
rect 18721 3349 18755 3383
rect 18889 3349 18923 3383
rect 22753 3349 22787 3383
rect 22845 3349 22879 3383
rect 22937 3349 22971 3383
rect 1961 3145 1995 3179
rect 11805 3145 11839 3179
rect 12081 3145 12115 3179
rect 15485 3145 15519 3179
rect 21281 3145 21315 3179
rect 21925 3145 21959 3179
rect 25053 3145 25087 3179
rect 13277 3077 13311 3111
rect 14933 3077 14967 3111
rect 15945 3077 15979 3111
rect 16129 3077 16163 3111
rect 16313 3077 16347 3111
rect 18153 3077 18187 3111
rect 19993 3077 20027 3111
rect 21097 3077 21131 3111
rect 22661 3077 22695 3111
rect 25237 3077 25271 3111
rect 28733 3077 28767 3111
rect 1593 3009 1627 3043
rect 1869 3009 1903 3043
rect 2145 3009 2179 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 13001 3009 13035 3043
rect 15025 3009 15059 3043
rect 15393 3009 15427 3043
rect 18429 3009 18463 3043
rect 20269 3009 20303 3043
rect 22017 3009 22051 3043
rect 22569 3009 22603 3043
rect 22753 3009 22787 3043
rect 22845 3009 22879 3043
rect 23029 3009 23063 3043
rect 23305 3009 23339 3043
rect 25329 3009 25363 3043
rect 28917 3009 28951 3043
rect 29285 3009 29319 3043
rect 16681 2941 16715 2975
rect 18521 2941 18555 2975
rect 20729 2941 20763 2975
rect 23581 2941 23615 2975
rect 1685 2873 1719 2907
rect 29101 2873 29135 2907
rect 14749 2805 14783 2839
rect 21097 2805 21131 2839
rect 23213 2805 23247 2839
rect 8309 2601 8343 2635
rect 9321 2601 9355 2635
rect 11897 2601 11931 2635
rect 15669 2601 15703 2635
rect 16221 2601 16255 2635
rect 17049 2601 17083 2635
rect 22845 2601 22879 2635
rect 23397 2601 23431 2635
rect 23581 2601 23615 2635
rect 23673 2601 23707 2635
rect 4997 2533 5031 2567
rect 20085 2533 20119 2567
rect 2329 2465 2363 2499
rect 5917 2465 5951 2499
rect 7481 2465 7515 2499
rect 24869 2465 24903 2499
rect 1777 2397 1811 2431
rect 2053 2397 2087 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 6193 2397 6227 2431
rect 7205 2397 7239 2431
rect 8125 2397 8159 2431
rect 9137 2397 9171 2431
rect 10425 2397 10459 2431
rect 10701 2397 10735 2431
rect 13001 2397 13035 2431
rect 13277 2397 13311 2431
rect 14565 2397 14599 2431
rect 16405 2397 16439 2431
rect 16957 2397 16991 2431
rect 17509 2397 17543 2431
rect 19441 2397 19475 2431
rect 20269 2397 20303 2431
rect 22661 2397 22695 2431
rect 23857 2397 23891 2431
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 28457 2397 28491 2431
rect 1501 2329 1535 2363
rect 4813 2329 4847 2363
rect 11805 2329 11839 2363
rect 14381 2329 14415 2363
rect 15761 2329 15795 2363
rect 18981 2329 19015 2363
rect 19349 2329 19383 2363
rect 23213 2329 23247 2363
rect 23413 2329 23447 2363
rect 26065 2329 26099 2363
rect 27353 2329 27387 2363
rect 28273 2329 28307 2363
rect 28641 2329 28675 2363
rect 29285 2329 29319 2363
rect 1593 2261 1627 2295
rect 1961 2261 1995 2295
rect 17739 2261 17773 2295
rect 18889 2261 18923 2295
rect 27261 2261 27295 2295
rect 28181 2261 28215 2295
rect 29193 2261 29227 2295
<< metal1 >>
rect 1104 30490 29716 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 29716 30490
rect 1104 30416 29716 30438
rect 1302 30268 1308 30320
rect 1360 30308 1366 30320
rect 2409 30311 2467 30317
rect 2409 30308 2421 30311
rect 1360 30280 2421 30308
rect 1360 30268 1366 30280
rect 2409 30277 2421 30280
rect 2455 30277 2467 30311
rect 2409 30271 2467 30277
rect 2590 30268 2596 30320
rect 2648 30308 2654 30320
rect 2777 30311 2835 30317
rect 2777 30308 2789 30311
rect 2648 30280 2789 30308
rect 2648 30268 2654 30280
rect 2777 30277 2789 30280
rect 2823 30277 2835 30311
rect 2777 30271 2835 30277
rect 8386 30268 8392 30320
rect 8444 30308 8450 30320
rect 8573 30311 8631 30317
rect 8573 30308 8585 30311
rect 8444 30280 8585 30308
rect 8444 30268 8450 30280
rect 8573 30277 8585 30280
rect 8619 30277 8631 30311
rect 8573 30271 8631 30277
rect 9674 30268 9680 30320
rect 9732 30308 9738 30320
rect 9861 30311 9919 30317
rect 9861 30308 9873 30311
rect 9732 30280 9873 30308
rect 9732 30268 9738 30280
rect 9861 30277 9873 30280
rect 9907 30277 9919 30311
rect 9861 30271 9919 30277
rect 15470 30268 15476 30320
rect 15528 30308 15534 30320
rect 15749 30311 15807 30317
rect 15749 30308 15761 30311
rect 15528 30280 15761 30308
rect 15528 30268 15534 30280
rect 15749 30277 15761 30280
rect 15795 30277 15807 30311
rect 15749 30271 15807 30277
rect 19334 30268 19340 30320
rect 19392 30308 19398 30320
rect 19613 30311 19671 30317
rect 19613 30308 19625 30311
rect 19392 30280 19625 30308
rect 19392 30268 19398 30280
rect 19613 30277 19625 30280
rect 19659 30277 19671 30311
rect 19613 30271 19671 30277
rect 20622 30268 20628 30320
rect 20680 30308 20686 30320
rect 20901 30311 20959 30317
rect 20901 30308 20913 30311
rect 20680 30280 20913 30308
rect 20680 30268 20686 30280
rect 20901 30277 20913 30280
rect 20947 30277 20959 30311
rect 20901 30271 20959 30277
rect 21910 30268 21916 30320
rect 21968 30308 21974 30320
rect 22097 30311 22155 30317
rect 22097 30308 22109 30311
rect 21968 30280 22109 30308
rect 21968 30268 21974 30280
rect 22097 30277 22109 30280
rect 22143 30277 22155 30311
rect 22097 30271 22155 30277
rect 25130 30268 25136 30320
rect 25188 30308 25194 30320
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 25188 30280 25421 30308
rect 25188 30268 25194 30280
rect 25409 30277 25421 30280
rect 25455 30277 25467 30311
rect 25409 30271 25467 30277
rect 27706 30268 27712 30320
rect 27764 30308 27770 30320
rect 28077 30311 28135 30317
rect 28077 30308 28089 30311
rect 27764 30280 28089 30308
rect 27764 30268 27770 30280
rect 28077 30277 28089 30280
rect 28123 30277 28135 30311
rect 30282 30308 30288 30320
rect 28077 30271 28135 30277
rect 28460 30280 30288 30308
rect 14 30200 20 30252
rect 72 30240 78 30252
rect 3145 30243 3203 30249
rect 72 30212 2774 30240
rect 72 30200 78 30212
rect 842 30132 848 30184
rect 900 30172 906 30184
rect 1397 30175 1455 30181
rect 1397 30172 1409 30175
rect 900 30144 1409 30172
rect 900 30132 906 30144
rect 1397 30141 1409 30144
rect 1443 30141 1455 30175
rect 1397 30135 1455 30141
rect 1673 30175 1731 30181
rect 1673 30141 1685 30175
rect 1719 30172 1731 30175
rect 1946 30172 1952 30184
rect 1719 30144 1952 30172
rect 1719 30141 1731 30144
rect 1673 30135 1731 30141
rect 1946 30132 1952 30144
rect 2004 30132 2010 30184
rect 2746 30172 2774 30212
rect 3145 30209 3157 30243
rect 3191 30209 3203 30243
rect 3145 30203 3203 30209
rect 3160 30172 3188 30203
rect 3878 30200 3884 30252
rect 3936 30240 3942 30252
rect 3973 30243 4031 30249
rect 3973 30240 3985 30243
rect 3936 30212 3985 30240
rect 3936 30200 3942 30212
rect 3973 30209 3985 30212
rect 4019 30209 4031 30243
rect 3973 30203 4031 30209
rect 5258 30200 5264 30252
rect 5316 30200 5322 30252
rect 7098 30200 7104 30252
rect 7156 30240 7162 30252
rect 7193 30243 7251 30249
rect 7193 30240 7205 30243
rect 7156 30212 7205 30240
rect 7156 30200 7162 30212
rect 7193 30209 7205 30212
rect 7239 30209 7251 30243
rect 7193 30203 7251 30209
rect 10962 30200 10968 30252
rect 11020 30240 11026 30252
rect 11057 30243 11115 30249
rect 11057 30240 11069 30243
rect 11020 30212 11069 30240
rect 11020 30200 11026 30212
rect 11057 30209 11069 30212
rect 11103 30209 11115 30243
rect 11057 30203 11115 30209
rect 12250 30200 12256 30252
rect 12308 30240 12314 30252
rect 12345 30243 12403 30249
rect 12345 30240 12357 30243
rect 12308 30212 12357 30240
rect 12308 30200 12314 30212
rect 12345 30209 12357 30212
rect 12391 30209 12403 30243
rect 12345 30203 12403 30209
rect 13538 30200 13544 30252
rect 13596 30240 13602 30252
rect 13817 30243 13875 30249
rect 13817 30240 13829 30243
rect 13596 30212 13829 30240
rect 13596 30200 13602 30212
rect 13817 30209 13829 30212
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 14826 30200 14832 30252
rect 14884 30240 14890 30252
rect 14921 30243 14979 30249
rect 14921 30240 14933 30243
rect 14884 30212 14933 30240
rect 14884 30200 14890 30212
rect 14921 30209 14933 30212
rect 14967 30209 14979 30243
rect 14921 30203 14979 30209
rect 16758 30200 16764 30252
rect 16816 30240 16822 30252
rect 16853 30243 16911 30249
rect 16853 30240 16865 30243
rect 16816 30212 16865 30240
rect 16816 30200 16822 30212
rect 16853 30209 16865 30212
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 18046 30200 18052 30252
rect 18104 30240 18110 30252
rect 18141 30243 18199 30249
rect 18141 30240 18153 30243
rect 18104 30212 18153 30240
rect 18104 30200 18110 30212
rect 18141 30209 18153 30212
rect 18187 30209 18199 30243
rect 18141 30203 18199 30209
rect 22554 30200 22560 30252
rect 22612 30240 22618 30252
rect 22649 30243 22707 30249
rect 22649 30240 22661 30243
rect 22612 30212 22661 30240
rect 22612 30200 22618 30212
rect 22649 30209 22661 30212
rect 22695 30209 22707 30243
rect 22649 30203 22707 30209
rect 23842 30200 23848 30252
rect 23900 30240 23906 30252
rect 23937 30243 23995 30249
rect 23937 30240 23949 30243
rect 23900 30212 23949 30240
rect 23900 30200 23906 30212
rect 23937 30209 23949 30212
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 28460 30249 28488 30280
rect 30282 30268 30288 30280
rect 30340 30268 30346 30320
rect 26973 30243 27031 30249
rect 26973 30240 26985 30243
rect 26476 30212 26985 30240
rect 26476 30200 26482 30212
rect 26973 30209 26985 30212
rect 27019 30209 27031 30243
rect 26973 30203 27031 30209
rect 28445 30243 28503 30249
rect 28445 30209 28457 30243
rect 28491 30209 28503 30243
rect 28445 30203 28503 30209
rect 29362 30200 29368 30252
rect 29420 30200 29426 30252
rect 11606 30172 11612 30184
rect 2746 30144 3188 30172
rect 7392 30144 11612 30172
rect 2593 30107 2651 30113
rect 2593 30073 2605 30107
rect 2639 30104 2651 30107
rect 2682 30104 2688 30116
rect 2639 30076 2688 30104
rect 2639 30073 2651 30076
rect 2593 30067 2651 30073
rect 2682 30064 2688 30076
rect 2740 30064 2746 30116
rect 2958 30064 2964 30116
rect 3016 30064 3022 30116
rect 3326 30064 3332 30116
rect 3384 30064 3390 30116
rect 7392 30113 7420 30144
rect 11606 30132 11612 30144
rect 11664 30132 11670 30184
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 17129 30175 17187 30181
rect 17129 30172 17141 30175
rect 16632 30144 17141 30172
rect 16632 30132 16638 30144
rect 17129 30141 17141 30144
rect 17175 30141 17187 30175
rect 17129 30135 17187 30141
rect 26510 30132 26516 30184
rect 26568 30172 26574 30184
rect 27249 30175 27307 30181
rect 27249 30172 27261 30175
rect 26568 30144 27261 30172
rect 26568 30132 26574 30144
rect 27249 30141 27261 30144
rect 27295 30141 27307 30175
rect 27249 30135 27307 30141
rect 29089 30175 29147 30181
rect 29089 30141 29101 30175
rect 29135 30172 29147 30175
rect 29730 30172 29736 30184
rect 29135 30144 29736 30172
rect 29135 30141 29147 30144
rect 29089 30135 29147 30141
rect 29730 30132 29736 30144
rect 29788 30132 29794 30184
rect 7377 30107 7435 30113
rect 7377 30073 7389 30107
rect 7423 30073 7435 30107
rect 7377 30067 7435 30073
rect 8757 30107 8815 30113
rect 8757 30073 8769 30107
rect 8803 30104 8815 30107
rect 9490 30104 9496 30116
rect 8803 30076 9496 30104
rect 8803 30073 8815 30076
rect 8757 30067 8815 30073
rect 9490 30064 9496 30076
rect 9548 30064 9554 30116
rect 10045 30107 10103 30113
rect 10045 30073 10057 30107
rect 10091 30104 10103 30107
rect 12066 30104 12072 30116
rect 10091 30076 12072 30104
rect 10091 30073 10103 30076
rect 10045 30067 10103 30073
rect 12066 30064 12072 30076
rect 12124 30064 12130 30116
rect 20714 30064 20720 30116
rect 20772 30064 20778 30116
rect 22281 30107 22339 30113
rect 22281 30073 22293 30107
rect 22327 30104 22339 30107
rect 22370 30104 22376 30116
rect 22327 30076 22376 30104
rect 22327 30073 22339 30076
rect 22281 30067 22339 30073
rect 22370 30064 22376 30076
rect 22428 30064 22434 30116
rect 27798 30064 27804 30116
rect 27856 30104 27862 30116
rect 27893 30107 27951 30113
rect 27893 30104 27905 30107
rect 27856 30076 27905 30104
rect 27856 30064 27862 30076
rect 27893 30073 27905 30076
rect 27939 30073 27951 30107
rect 27893 30067 27951 30073
rect 4157 30039 4215 30045
rect 4157 30005 4169 30039
rect 4203 30036 4215 30039
rect 5258 30036 5264 30048
rect 4203 30008 5264 30036
rect 4203 30005 4215 30008
rect 4157 29999 4215 30005
rect 5258 29996 5264 30008
rect 5316 29996 5322 30048
rect 5442 29996 5448 30048
rect 5500 29996 5506 30048
rect 11241 30039 11299 30045
rect 11241 30005 11253 30039
rect 11287 30036 11299 30039
rect 12158 30036 12164 30048
rect 11287 30008 12164 30036
rect 11287 30005 11299 30008
rect 11241 29999 11299 30005
rect 12158 29996 12164 30008
rect 12216 29996 12222 30048
rect 12526 29996 12532 30048
rect 12584 29996 12590 30048
rect 13538 29996 13544 30048
rect 13596 30036 13602 30048
rect 13633 30039 13691 30045
rect 13633 30036 13645 30039
rect 13596 30008 13645 30036
rect 13596 29996 13602 30008
rect 13633 30005 13645 30008
rect 13679 30005 13691 30039
rect 13633 29999 13691 30005
rect 14918 29996 14924 30048
rect 14976 30036 14982 30048
rect 15105 30039 15163 30045
rect 15105 30036 15117 30039
rect 14976 30008 15117 30036
rect 14976 29996 14982 30008
rect 15105 30005 15117 30008
rect 15151 30005 15163 30039
rect 15105 29999 15163 30005
rect 15654 29996 15660 30048
rect 15712 29996 15718 30048
rect 18322 29996 18328 30048
rect 18380 29996 18386 30048
rect 19518 29996 19524 30048
rect 19576 29996 19582 30048
rect 22833 30039 22891 30045
rect 22833 30005 22845 30039
rect 22879 30036 22891 30039
rect 23934 30036 23940 30048
rect 22879 30008 23940 30036
rect 22879 30005 22891 30008
rect 22833 29999 22891 30005
rect 23934 29996 23940 30008
rect 23992 29996 23998 30048
rect 24118 29996 24124 30048
rect 24176 29996 24182 30048
rect 25317 30039 25375 30045
rect 25317 30005 25329 30039
rect 25363 30036 25375 30039
rect 26142 30036 26148 30048
rect 25363 30008 26148 30036
rect 25363 30005 25375 30008
rect 25317 29999 25375 30005
rect 26142 29996 26148 30008
rect 26200 29996 26206 30048
rect 28074 29996 28080 30048
rect 28132 30036 28138 30048
rect 28261 30039 28319 30045
rect 28261 30036 28273 30039
rect 28132 30008 28273 30036
rect 28132 29996 28138 30008
rect 28261 30005 28273 30008
rect 28307 30005 28319 30039
rect 28261 29999 28319 30005
rect 1104 29946 29716 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 29716 29946
rect 1104 29872 29716 29894
rect 934 29656 940 29708
rect 992 29696 998 29708
rect 1397 29699 1455 29705
rect 1397 29696 1409 29699
rect 992 29668 1409 29696
rect 992 29656 998 29668
rect 1397 29665 1409 29668
rect 1443 29665 1455 29699
rect 1397 29659 1455 29665
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 9214 29628 9220 29640
rect 1719 29600 9220 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 13538 29588 13544 29640
rect 13596 29588 13602 29640
rect 28534 29588 28540 29640
rect 28592 29588 28598 29640
rect 28902 29588 28908 29640
rect 28960 29588 28966 29640
rect 28994 29588 29000 29640
rect 29052 29628 29058 29640
rect 29273 29631 29331 29637
rect 29273 29628 29285 29631
rect 29052 29600 29285 29628
rect 29052 29588 29058 29600
rect 29273 29597 29285 29600
rect 29319 29597 29331 29631
rect 29273 29591 29331 29597
rect 1210 29520 1216 29572
rect 1268 29560 1274 29572
rect 2409 29563 2467 29569
rect 2409 29560 2421 29563
rect 1268 29532 2421 29560
rect 1268 29520 1274 29532
rect 2409 29529 2421 29532
rect 2455 29529 2467 29563
rect 2409 29523 2467 29529
rect 2590 29520 2596 29572
rect 2648 29520 2654 29572
rect 28350 29520 28356 29572
rect 28408 29520 28414 29572
rect 28626 29520 28632 29572
rect 28684 29560 28690 29572
rect 28721 29563 28779 29569
rect 28721 29560 28733 29563
rect 28684 29532 28733 29560
rect 28684 29520 28690 29532
rect 28721 29529 28733 29532
rect 28767 29529 28779 29563
rect 28721 29523 28779 29529
rect 13078 29452 13084 29504
rect 13136 29492 13142 29504
rect 13449 29495 13507 29501
rect 13449 29492 13461 29495
rect 13136 29464 13461 29492
rect 13136 29452 13142 29464
rect 13449 29461 13461 29464
rect 13495 29461 13507 29495
rect 13449 29455 13507 29461
rect 29181 29495 29239 29501
rect 29181 29461 29193 29495
rect 29227 29492 29239 29495
rect 29454 29492 29460 29504
rect 29227 29464 29460 29492
rect 29227 29461 29239 29464
rect 29181 29455 29239 29461
rect 29454 29452 29460 29464
rect 29512 29452 29518 29504
rect 1104 29402 29716 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 29716 29402
rect 1104 29328 29716 29350
rect 17862 29248 17868 29300
rect 17920 29288 17926 29300
rect 19521 29291 19579 29297
rect 19521 29288 19533 29291
rect 17920 29260 19533 29288
rect 17920 29248 17926 29260
rect 19521 29257 19533 29260
rect 19567 29257 19579 29291
rect 19521 29251 19579 29257
rect 15746 29180 15752 29232
rect 15804 29180 15810 29232
rect 18782 29180 18788 29232
rect 18840 29180 18846 29232
rect 1394 29112 1400 29164
rect 1452 29112 1458 29164
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29152 11207 29155
rect 12434 29152 12440 29164
rect 11195 29124 12440 29152
rect 11195 29121 11207 29124
rect 11149 29115 11207 29121
rect 12434 29112 12440 29124
rect 12492 29152 12498 29164
rect 13630 29152 13636 29164
rect 12492 29124 13636 29152
rect 12492 29112 12498 29124
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 21082 29112 21088 29164
rect 21140 29152 21146 29164
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 21140 29124 23121 29152
rect 21140 29112 21146 29124
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 23109 29115 23167 29121
rect 29270 29112 29276 29164
rect 29328 29112 29334 29164
rect 3145 29087 3203 29093
rect 3145 29053 3157 29087
rect 3191 29084 3203 29087
rect 4706 29084 4712 29096
rect 3191 29056 4712 29084
rect 3191 29053 3203 29056
rect 3145 29047 3203 29053
rect 4706 29044 4712 29056
rect 4764 29044 4770 29096
rect 12618 29044 12624 29096
rect 12676 29084 12682 29096
rect 14461 29087 14519 29093
rect 14461 29084 14473 29087
rect 12676 29056 14473 29084
rect 12676 29044 12682 29056
rect 14461 29053 14473 29056
rect 14507 29053 14519 29087
rect 14461 29047 14519 29053
rect 15470 29044 15476 29096
rect 15528 29084 15534 29096
rect 16485 29087 16543 29093
rect 16485 29084 16497 29087
rect 15528 29056 16497 29084
rect 15528 29044 15534 29056
rect 16485 29053 16497 29056
rect 16531 29053 16543 29087
rect 16485 29047 16543 29053
rect 17773 29087 17831 29093
rect 17773 29053 17785 29087
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 11146 28976 11152 29028
rect 11204 29016 11210 29028
rect 11241 29019 11299 29025
rect 11241 29016 11253 29019
rect 11204 28988 11253 29016
rect 11204 28976 11210 28988
rect 11241 28985 11253 28988
rect 11287 28985 11299 29019
rect 17788 29016 17816 29047
rect 18046 29044 18052 29096
rect 18104 29044 18110 29096
rect 23201 29019 23259 29025
rect 17788 28988 17908 29016
rect 11241 28979 11299 28985
rect 14550 28908 14556 28960
rect 14608 28948 14614 28960
rect 14718 28951 14776 28957
rect 14718 28948 14730 28951
rect 14608 28920 14730 28948
rect 14608 28908 14614 28920
rect 14718 28917 14730 28920
rect 14764 28917 14776 28951
rect 17880 28948 17908 28988
rect 23201 28985 23213 29019
rect 23247 29016 23259 29019
rect 23474 29016 23480 29028
rect 23247 28988 23480 29016
rect 23247 28985 23259 28988
rect 23201 28979 23259 28985
rect 23474 28976 23480 28988
rect 23532 28976 23538 29028
rect 29089 29019 29147 29025
rect 29089 28985 29101 29019
rect 29135 29016 29147 29019
rect 29178 29016 29184 29028
rect 29135 28988 29184 29016
rect 29135 28985 29147 28988
rect 29089 28979 29147 28985
rect 29178 28976 29184 28988
rect 29236 28976 29242 29028
rect 18506 28948 18512 28960
rect 17880 28920 18512 28948
rect 14718 28911 14776 28917
rect 18506 28908 18512 28920
rect 18564 28908 18570 28960
rect 1104 28858 29716 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 29716 28858
rect 1104 28784 29716 28806
rect 5258 28704 5264 28756
rect 5316 28744 5322 28756
rect 9306 28744 9312 28756
rect 5316 28716 9312 28744
rect 5316 28704 5322 28716
rect 9306 28704 9312 28716
rect 9364 28704 9370 28756
rect 15657 28747 15715 28753
rect 15657 28713 15669 28747
rect 15703 28744 15715 28747
rect 15746 28744 15752 28756
rect 15703 28716 15752 28744
rect 15703 28713 15715 28716
rect 15657 28707 15715 28713
rect 15746 28704 15752 28716
rect 15804 28704 15810 28756
rect 18782 28704 18788 28756
rect 18840 28744 18846 28756
rect 18877 28747 18935 28753
rect 18877 28744 18889 28747
rect 18840 28716 18889 28744
rect 18840 28704 18846 28716
rect 18877 28713 18889 28716
rect 18923 28713 18935 28747
rect 18877 28707 18935 28713
rect 8113 28679 8171 28685
rect 8113 28676 8125 28679
rect 7484 28648 8125 28676
rect 7282 28500 7288 28552
rect 7340 28500 7346 28552
rect 7484 28549 7512 28648
rect 8113 28645 8125 28648
rect 8159 28645 8171 28679
rect 8113 28639 8171 28645
rect 25314 28636 25320 28688
rect 25372 28676 25378 28688
rect 25777 28679 25835 28685
rect 25777 28676 25789 28679
rect 25372 28648 25789 28676
rect 25372 28636 25378 28648
rect 25777 28645 25789 28648
rect 25823 28645 25835 28679
rect 25777 28639 25835 28645
rect 10410 28568 10416 28620
rect 10468 28608 10474 28620
rect 12161 28611 12219 28617
rect 12161 28608 12173 28611
rect 10468 28580 12173 28608
rect 10468 28568 10474 28580
rect 12161 28577 12173 28580
rect 12207 28577 12219 28611
rect 12161 28571 12219 28577
rect 17221 28611 17279 28617
rect 17221 28577 17233 28611
rect 17267 28608 17279 28611
rect 17267 28580 17816 28608
rect 17267 28577 17279 28580
rect 17221 28571 17279 28577
rect 7469 28543 7527 28549
rect 7469 28509 7481 28543
rect 7515 28509 7527 28543
rect 7469 28503 7527 28509
rect 7558 28500 7564 28552
rect 7616 28500 7622 28552
rect 7653 28543 7711 28549
rect 7653 28509 7665 28543
rect 7699 28509 7711 28543
rect 7653 28503 7711 28509
rect 7466 28364 7472 28416
rect 7524 28404 7530 28416
rect 7668 28404 7696 28503
rect 8202 28500 8208 28552
rect 8260 28500 8266 28552
rect 9122 28500 9128 28552
rect 9180 28500 9186 28552
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28509 10195 28543
rect 10137 28503 10195 28509
rect 10152 28472 10180 28503
rect 12342 28500 12348 28552
rect 12400 28540 12406 28552
rect 12437 28543 12495 28549
rect 12437 28540 12449 28543
rect 12400 28512 12449 28540
rect 12400 28500 12406 28512
rect 12437 28509 12449 28512
rect 12483 28509 12495 28543
rect 12437 28503 12495 28509
rect 12621 28543 12679 28549
rect 12621 28509 12633 28543
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 10413 28475 10471 28481
rect 10152 28444 10272 28472
rect 7524 28376 7696 28404
rect 7929 28407 7987 28413
rect 7524 28364 7530 28376
rect 7929 28373 7941 28407
rect 7975 28404 7987 28407
rect 8018 28404 8024 28416
rect 7975 28376 8024 28404
rect 7975 28373 7987 28376
rect 7929 28367 7987 28373
rect 8018 28364 8024 28376
rect 8076 28364 8082 28416
rect 9030 28364 9036 28416
rect 9088 28364 9094 28416
rect 10244 28404 10272 28444
rect 10413 28441 10425 28475
rect 10459 28472 10471 28475
rect 10502 28472 10508 28484
rect 10459 28444 10508 28472
rect 10459 28441 10471 28444
rect 10413 28435 10471 28441
rect 10502 28432 10508 28444
rect 10560 28432 10566 28484
rect 11146 28432 11152 28484
rect 11204 28432 11210 28484
rect 12636 28472 12664 28503
rect 12710 28500 12716 28552
rect 12768 28500 12774 28552
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28540 12863 28543
rect 13170 28540 13176 28552
rect 12851 28512 13176 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 13170 28500 13176 28512
rect 13228 28500 13234 28552
rect 13630 28500 13636 28552
rect 13688 28540 13694 28552
rect 15749 28543 15807 28549
rect 15749 28540 15761 28543
rect 13688 28512 15761 28540
rect 13688 28500 13694 28512
rect 15749 28509 15761 28512
rect 15795 28540 15807 28543
rect 16942 28540 16948 28552
rect 15795 28512 16948 28540
rect 15795 28509 15807 28512
rect 15749 28503 15807 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17402 28500 17408 28552
rect 17460 28540 17466 28552
rect 17681 28543 17739 28549
rect 17681 28540 17693 28543
rect 17460 28512 17693 28540
rect 17460 28500 17466 28512
rect 17681 28509 17693 28512
rect 17727 28509 17739 28543
rect 17788 28540 17816 28580
rect 18506 28568 18512 28620
rect 18564 28608 18570 28620
rect 19978 28608 19984 28620
rect 18564 28580 19984 28608
rect 18564 28568 18570 28580
rect 19978 28568 19984 28580
rect 20036 28608 20042 28620
rect 22189 28611 22247 28617
rect 22189 28608 22201 28611
rect 20036 28580 22201 28608
rect 20036 28568 20042 28580
rect 22189 28577 22201 28580
rect 22235 28577 22247 28611
rect 22189 28571 22247 28577
rect 22465 28611 22523 28617
rect 22465 28577 22477 28611
rect 22511 28608 22523 28611
rect 24121 28611 24179 28617
rect 24121 28608 24133 28611
rect 22511 28580 24133 28608
rect 22511 28577 22523 28580
rect 22465 28571 22523 28577
rect 24121 28577 24133 28580
rect 24167 28577 24179 28611
rect 24121 28571 24179 28577
rect 17862 28540 17868 28552
rect 17920 28549 17926 28552
rect 17788 28512 17868 28540
rect 17681 28503 17739 28509
rect 17862 28500 17868 28512
rect 17920 28540 17931 28549
rect 18230 28540 18236 28552
rect 17920 28512 18236 28540
rect 17920 28503 17931 28512
rect 17920 28500 17926 28503
rect 18230 28500 18236 28512
rect 18288 28500 18294 28552
rect 18785 28543 18843 28549
rect 18785 28509 18797 28543
rect 18831 28509 18843 28543
rect 18785 28503 18843 28509
rect 13998 28472 14004 28484
rect 12636 28444 14004 28472
rect 13998 28432 14004 28444
rect 14056 28432 14062 28484
rect 16960 28472 16988 28500
rect 18800 28472 18828 28503
rect 24026 28500 24032 28552
rect 24084 28500 24090 28552
rect 24213 28543 24271 28549
rect 24213 28509 24225 28543
rect 24259 28540 24271 28543
rect 24486 28540 24492 28552
rect 24259 28512 24492 28540
rect 24259 28509 24271 28512
rect 24213 28503 24271 28509
rect 24486 28500 24492 28512
rect 24544 28500 24550 28552
rect 25498 28500 25504 28552
rect 25556 28500 25562 28552
rect 27062 28500 27068 28552
rect 27120 28500 27126 28552
rect 29086 28500 29092 28552
rect 29144 28500 29150 28552
rect 16960 28444 18828 28472
rect 11330 28404 11336 28416
rect 10244 28376 11336 28404
rect 11330 28364 11336 28376
rect 11388 28364 11394 28416
rect 12894 28364 12900 28416
rect 12952 28404 12958 28416
rect 13081 28407 13139 28413
rect 13081 28404 13093 28407
rect 12952 28376 13093 28404
rect 12952 28364 12958 28376
rect 13081 28373 13093 28376
rect 13127 28373 13139 28407
rect 13081 28367 13139 28373
rect 13630 28364 13636 28416
rect 13688 28404 13694 28416
rect 13725 28407 13783 28413
rect 13725 28404 13737 28407
rect 13688 28376 13737 28404
rect 13688 28364 13694 28376
rect 13725 28373 13737 28376
rect 13771 28373 13783 28407
rect 13725 28367 13783 28373
rect 17586 28364 17592 28416
rect 17644 28364 17650 28416
rect 17954 28364 17960 28416
rect 18012 28404 18018 28416
rect 18049 28407 18107 28413
rect 18049 28404 18061 28407
rect 18012 28376 18061 28404
rect 18012 28364 18018 28376
rect 18049 28373 18061 28376
rect 18095 28373 18107 28407
rect 18800 28404 18828 28444
rect 20254 28432 20260 28484
rect 20312 28432 20318 28484
rect 21266 28432 21272 28484
rect 21324 28432 21330 28484
rect 22002 28432 22008 28484
rect 22060 28432 22066 28484
rect 23474 28432 23480 28484
rect 23532 28432 23538 28484
rect 25774 28432 25780 28484
rect 25832 28432 25838 28484
rect 27338 28432 27344 28484
rect 27396 28432 27402 28484
rect 28997 28475 29055 28481
rect 28997 28472 29009 28475
rect 28566 28444 29009 28472
rect 28997 28441 29009 28444
rect 29043 28441 29055 28475
rect 28997 28435 29055 28441
rect 21082 28404 21088 28416
rect 18800 28376 21088 28404
rect 18049 28367 18107 28373
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 23937 28407 23995 28413
rect 23937 28373 23949 28407
rect 23983 28404 23995 28407
rect 24210 28404 24216 28416
rect 23983 28376 24216 28404
rect 23983 28373 23995 28376
rect 23937 28367 23995 28373
rect 24210 28364 24216 28376
rect 24268 28364 24274 28416
rect 25593 28407 25651 28413
rect 25593 28373 25605 28407
rect 25639 28404 25651 28407
rect 25958 28404 25964 28416
rect 25639 28376 25964 28404
rect 25639 28373 25651 28376
rect 25593 28367 25651 28373
rect 25958 28364 25964 28376
rect 26016 28404 26022 28416
rect 27154 28404 27160 28416
rect 26016 28376 27160 28404
rect 26016 28364 26022 28376
rect 27154 28364 27160 28376
rect 27212 28404 27218 28416
rect 28813 28407 28871 28413
rect 28813 28404 28825 28407
rect 27212 28376 28825 28404
rect 27212 28364 27218 28376
rect 28813 28373 28825 28376
rect 28859 28373 28871 28407
rect 28813 28367 28871 28373
rect 1104 28314 29716 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 29716 28314
rect 1104 28240 29716 28262
rect 7282 28160 7288 28212
rect 7340 28200 7346 28212
rect 7340 28172 9904 28200
rect 7340 28160 7346 28172
rect 5828 28104 7420 28132
rect 4706 28024 4712 28076
rect 4764 28064 4770 28076
rect 5828 28073 5856 28104
rect 5813 28067 5871 28073
rect 5813 28064 5825 28067
rect 4764 28036 5825 28064
rect 4764 28024 4770 28036
rect 5813 28033 5825 28036
rect 5859 28033 5871 28067
rect 5813 28027 5871 28033
rect 5902 28024 5908 28076
rect 5960 28064 5966 28076
rect 6365 28067 6423 28073
rect 6365 28064 6377 28067
rect 5960 28036 6377 28064
rect 5960 28024 5966 28036
rect 6365 28033 6377 28036
rect 6411 28033 6423 28067
rect 6365 28027 6423 28033
rect 6380 27996 6408 28027
rect 6546 28024 6552 28076
rect 6604 28024 6610 28076
rect 7098 27996 7104 28008
rect 6380 27968 7104 27996
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 5810 27820 5816 27872
rect 5868 27860 5874 27872
rect 5905 27863 5963 27869
rect 5905 27860 5917 27863
rect 5868 27832 5917 27860
rect 5868 27820 5874 27832
rect 5905 27829 5917 27832
rect 5951 27829 5963 27863
rect 5905 27823 5963 27829
rect 6454 27820 6460 27872
rect 6512 27820 6518 27872
rect 7392 27860 7420 28104
rect 8018 28092 8024 28144
rect 8076 28092 8082 28144
rect 9030 28092 9036 28144
rect 9088 28092 9094 28144
rect 9876 28073 9904 28172
rect 10502 28160 10508 28212
rect 10560 28160 10566 28212
rect 10686 28160 10692 28212
rect 10744 28200 10750 28212
rect 11057 28203 11115 28209
rect 11057 28200 11069 28203
rect 10744 28172 11069 28200
rect 10744 28160 10750 28172
rect 11057 28169 11069 28172
rect 11103 28200 11115 28203
rect 12710 28200 12716 28212
rect 11103 28172 12716 28200
rect 11103 28169 11115 28172
rect 11057 28163 11115 28169
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 13170 28160 13176 28212
rect 13228 28200 13234 28212
rect 13906 28200 13912 28212
rect 13228 28172 13912 28200
rect 13228 28160 13234 28172
rect 13906 28160 13912 28172
rect 13964 28200 13970 28212
rect 14369 28203 14427 28209
rect 14369 28200 14381 28203
rect 13964 28172 14381 28200
rect 13964 28160 13970 28172
rect 14369 28169 14381 28172
rect 14415 28169 14427 28203
rect 14369 28163 14427 28169
rect 14550 28160 14556 28212
rect 14608 28160 14614 28212
rect 14826 28160 14832 28212
rect 14884 28200 14890 28212
rect 15489 28203 15547 28209
rect 15489 28200 15501 28203
rect 14884 28172 15501 28200
rect 14884 28160 14890 28172
rect 15489 28169 15501 28172
rect 15535 28169 15547 28203
rect 15489 28163 15547 28169
rect 15657 28203 15715 28209
rect 15657 28169 15669 28203
rect 15703 28200 15715 28203
rect 17402 28200 17408 28212
rect 15703 28172 17408 28200
rect 15703 28169 15715 28172
rect 15657 28163 15715 28169
rect 10704 28104 11008 28132
rect 9861 28067 9919 28073
rect 9861 28033 9873 28067
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 7742 27956 7748 28008
rect 7800 27956 7806 28008
rect 9769 27999 9827 28005
rect 9769 27996 9781 27999
rect 7852 27968 9781 27996
rect 7466 27888 7472 27940
rect 7524 27928 7530 27940
rect 7852 27928 7880 27968
rect 9769 27965 9781 27968
rect 9815 27965 9827 27999
rect 9769 27959 9827 27965
rect 7524 27900 7880 27928
rect 9876 27928 9904 28027
rect 10042 28024 10048 28076
rect 10100 28024 10106 28076
rect 10134 28024 10140 28076
rect 10192 28024 10198 28076
rect 10226 28024 10232 28076
rect 10284 28024 10290 28076
rect 10704 28073 10732 28104
rect 10980 28073 11008 28104
rect 12894 28092 12900 28144
rect 12952 28092 12958 28144
rect 13630 28092 13636 28144
rect 13688 28092 13694 28144
rect 14734 28092 14740 28144
rect 14792 28092 14798 28144
rect 15286 28092 15292 28144
rect 15344 28092 15350 28144
rect 10689 28067 10747 28073
rect 10689 28033 10701 28067
rect 10735 28033 10747 28067
rect 10689 28027 10747 28033
rect 10873 28067 10931 28073
rect 10873 28033 10885 28067
rect 10919 28033 10931 28067
rect 10873 28027 10931 28033
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 10060 27996 10088 28024
rect 10704 27996 10732 28027
rect 10060 27968 10732 27996
rect 10888 27996 10916 28027
rect 11146 28024 11152 28076
rect 11204 28024 11210 28076
rect 11330 28024 11336 28076
rect 11388 28064 11394 28076
rect 12618 28064 12624 28076
rect 11388 28036 12624 28064
rect 11388 28024 11394 28036
rect 12618 28024 12624 28036
rect 12676 28024 12682 28076
rect 15764 28073 15792 28172
rect 17402 28160 17408 28172
rect 17460 28160 17466 28212
rect 17586 28160 17592 28212
rect 17644 28200 17650 28212
rect 19061 28203 19119 28209
rect 17644 28172 18920 28200
rect 17644 28160 17650 28172
rect 16114 28092 16120 28144
rect 16172 28092 16178 28144
rect 18892 28132 18920 28172
rect 19061 28169 19073 28203
rect 19107 28200 19119 28203
rect 19242 28200 19248 28212
rect 19107 28172 19248 28200
rect 19107 28169 19119 28172
rect 19061 28163 19119 28169
rect 19242 28160 19248 28172
rect 19300 28200 19306 28212
rect 19813 28203 19871 28209
rect 19813 28200 19825 28203
rect 19300 28172 19825 28200
rect 19300 28160 19306 28172
rect 19813 28169 19825 28172
rect 19859 28169 19871 28203
rect 19813 28163 19871 28169
rect 19981 28203 20039 28209
rect 19981 28169 19993 28203
rect 20027 28200 20039 28203
rect 20254 28200 20260 28212
rect 20027 28172 20260 28200
rect 20027 28169 20039 28172
rect 19981 28163 20039 28169
rect 20254 28160 20260 28172
rect 20312 28160 20318 28212
rect 21177 28203 21235 28209
rect 21177 28169 21189 28203
rect 21223 28200 21235 28203
rect 21266 28200 21272 28212
rect 21223 28172 21272 28200
rect 21223 28169 21235 28172
rect 21177 28163 21235 28169
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 24486 28160 24492 28212
rect 24544 28160 24550 28212
rect 19153 28135 19211 28141
rect 19153 28132 19165 28135
rect 18892 28104 19165 28132
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 17126 28024 17132 28076
rect 17184 28024 17190 28076
rect 18506 28024 18512 28076
rect 18564 28024 18570 28076
rect 18892 28073 18920 28104
rect 19153 28101 19165 28104
rect 19199 28101 19211 28135
rect 19153 28095 19211 28101
rect 19426 28092 19432 28144
rect 19484 28132 19490 28144
rect 19613 28135 19671 28141
rect 19613 28132 19625 28135
rect 19484 28104 19625 28132
rect 19484 28092 19490 28104
rect 19613 28101 19625 28104
rect 19659 28101 19671 28135
rect 22002 28132 22008 28144
rect 19613 28095 19671 28101
rect 21192 28104 22008 28132
rect 18877 28067 18935 28073
rect 18877 28033 18889 28067
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 18966 28024 18972 28076
rect 19024 28064 19030 28076
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 19024 28036 19073 28064
rect 19024 28024 19030 28036
rect 19061 28033 19073 28036
rect 19107 28064 19119 28067
rect 19337 28067 19395 28073
rect 19337 28064 19349 28067
rect 19107 28036 19349 28064
rect 19107 28033 19119 28036
rect 19061 28027 19119 28033
rect 19337 28033 19349 28036
rect 19383 28064 19395 28067
rect 21192 28064 21220 28104
rect 22002 28092 22008 28104
rect 22060 28092 22066 28144
rect 25130 28132 25136 28144
rect 24136 28104 25136 28132
rect 19383 28036 21220 28064
rect 21269 28067 21327 28073
rect 19383 28033 19395 28036
rect 19337 28027 19395 28033
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 11164 27996 11192 28024
rect 18233 27999 18291 28005
rect 18233 27996 18245 27999
rect 10888 27968 11192 27996
rect 16316 27968 18245 27996
rect 11054 27928 11060 27940
rect 9876 27900 11060 27928
rect 7524 27888 7530 27900
rect 11054 27888 11060 27900
rect 11112 27928 11118 27940
rect 12342 27928 12348 27940
rect 11112 27900 12348 27928
rect 11112 27888 11118 27900
rect 12342 27888 12348 27900
rect 12400 27928 12406 27940
rect 12400 27888 12434 27928
rect 14182 27888 14188 27940
rect 14240 27928 14246 27940
rect 15010 27928 15016 27940
rect 14240 27900 15016 27928
rect 14240 27888 14246 27900
rect 15010 27888 15016 27900
rect 15068 27928 15074 27940
rect 16316 27937 16344 27968
rect 18233 27965 18245 27968
rect 18279 27965 18291 27999
rect 18233 27959 18291 27965
rect 21082 27956 21088 28008
rect 21140 27996 21146 28008
rect 21284 27996 21312 28027
rect 23474 28024 23480 28076
rect 23532 28024 23538 28076
rect 24136 28073 24164 28104
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28033 24179 28067
rect 24121 28027 24179 28033
rect 24210 28024 24216 28076
rect 24268 28064 24274 28076
rect 24596 28073 24624 28104
rect 25130 28092 25136 28104
rect 25188 28092 25194 28144
rect 26697 28135 26755 28141
rect 26697 28132 26709 28135
rect 26266 28104 26709 28132
rect 26697 28101 26709 28104
rect 26743 28101 26755 28135
rect 29086 28132 29092 28144
rect 26697 28095 26755 28101
rect 26804 28104 29092 28132
rect 26804 28073 26832 28104
rect 29086 28092 29092 28104
rect 29144 28092 29150 28144
rect 24397 28067 24455 28073
rect 24397 28064 24409 28067
rect 24268 28036 24409 28064
rect 24268 28024 24274 28036
rect 24397 28033 24409 28036
rect 24443 28033 24455 28067
rect 24397 28027 24455 28033
rect 24581 28067 24639 28073
rect 24581 28033 24593 28067
rect 24627 28033 24639 28067
rect 24581 28027 24639 28033
rect 26789 28067 26847 28073
rect 26789 28033 26801 28067
rect 26835 28033 26847 28067
rect 26789 28027 26847 28033
rect 27154 28024 27160 28076
rect 27212 28024 27218 28076
rect 21140 27968 21312 27996
rect 23569 27999 23627 28005
rect 21140 27956 21146 27968
rect 23569 27965 23581 27999
rect 23615 27996 23627 27999
rect 23658 27996 23664 28008
rect 23615 27968 23664 27996
rect 23615 27965 23627 27968
rect 23569 27959 23627 27965
rect 23658 27956 23664 27968
rect 23716 27996 23722 28008
rect 23937 27999 23995 28005
rect 23937 27996 23949 27999
rect 23716 27968 23949 27996
rect 23716 27956 23722 27968
rect 23937 27965 23949 27968
rect 23983 27996 23995 27999
rect 24026 27996 24032 28008
rect 23983 27968 24032 27996
rect 23983 27965 23995 27968
rect 23937 27959 23995 27965
rect 24026 27956 24032 27968
rect 24084 27956 24090 28008
rect 24762 27956 24768 28008
rect 24820 27956 24826 28008
rect 25038 27956 25044 28008
rect 25096 27956 25102 28008
rect 25774 27956 25780 28008
rect 25832 27996 25838 28008
rect 26513 27999 26571 28005
rect 26513 27996 26525 27999
rect 25832 27968 26525 27996
rect 25832 27956 25838 27968
rect 26513 27965 26525 27968
rect 26559 27965 26571 27999
rect 26513 27959 26571 27965
rect 27065 27999 27123 28005
rect 27065 27965 27077 27999
rect 27111 27965 27123 27999
rect 27065 27959 27123 27965
rect 15105 27931 15163 27937
rect 15105 27928 15117 27931
rect 15068 27900 15117 27928
rect 15068 27888 15074 27900
rect 15105 27897 15117 27900
rect 15151 27897 15163 27931
rect 16301 27931 16359 27937
rect 15105 27891 15163 27897
rect 15396 27900 16160 27928
rect 9122 27860 9128 27872
rect 7392 27832 9128 27860
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 10778 27820 10784 27872
rect 10836 27820 10842 27872
rect 12406 27860 12434 27888
rect 14642 27860 14648 27872
rect 12406 27832 14648 27860
rect 14642 27820 14648 27832
rect 14700 27860 14706 27872
rect 14737 27863 14795 27869
rect 14737 27860 14749 27863
rect 14700 27832 14749 27860
rect 14700 27820 14706 27832
rect 14737 27829 14749 27832
rect 14783 27860 14795 27863
rect 15396 27860 15424 27900
rect 14783 27832 15424 27860
rect 14783 27829 14795 27832
rect 14737 27823 14795 27829
rect 15470 27820 15476 27872
rect 15528 27820 15534 27872
rect 16132 27869 16160 27900
rect 16301 27897 16313 27931
rect 16347 27897 16359 27931
rect 16301 27891 16359 27897
rect 16117 27863 16175 27869
rect 16117 27829 16129 27863
rect 16163 27860 16175 27863
rect 16390 27860 16396 27872
rect 16163 27832 16396 27860
rect 16163 27829 16175 27832
rect 16117 27823 16175 27829
rect 16390 27820 16396 27832
rect 16448 27820 16454 27872
rect 16758 27820 16764 27872
rect 16816 27820 16822 27872
rect 17862 27820 17868 27872
rect 17920 27860 17926 27872
rect 19426 27860 19432 27872
rect 17920 27832 19432 27860
rect 17920 27820 17926 27832
rect 19426 27820 19432 27832
rect 19484 27820 19490 27872
rect 19521 27863 19579 27869
rect 19521 27829 19533 27863
rect 19567 27860 19579 27863
rect 19797 27863 19855 27869
rect 19797 27860 19809 27863
rect 19567 27832 19809 27860
rect 19567 27829 19579 27832
rect 19521 27823 19579 27829
rect 19797 27829 19809 27832
rect 19843 27829 19855 27863
rect 19797 27823 19855 27829
rect 23842 27820 23848 27872
rect 23900 27820 23906 27872
rect 25498 27820 25504 27872
rect 25556 27860 25562 27872
rect 27080 27860 27108 27959
rect 27338 27956 27344 28008
rect 27396 27996 27402 28008
rect 27525 27999 27583 28005
rect 27525 27996 27537 27999
rect 27396 27968 27537 27996
rect 27396 27956 27402 27968
rect 27525 27965 27537 27968
rect 27571 27965 27583 27999
rect 27525 27959 27583 27965
rect 25556 27832 27108 27860
rect 25556 27820 25562 27832
rect 1104 27770 29716 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 29716 27770
rect 1104 27696 29716 27718
rect 7285 27659 7343 27665
rect 7285 27625 7297 27659
rect 7331 27656 7343 27659
rect 8297 27659 8355 27665
rect 8297 27656 8309 27659
rect 7331 27628 8309 27656
rect 7331 27625 7343 27628
rect 7285 27619 7343 27625
rect 8297 27625 8309 27628
rect 8343 27625 8355 27659
rect 8297 27619 8355 27625
rect 9953 27659 10011 27665
rect 9953 27625 9965 27659
rect 9999 27656 10011 27659
rect 10042 27656 10048 27668
rect 9999 27628 10048 27656
rect 9999 27625 10011 27628
rect 9953 27619 10011 27625
rect 10042 27616 10048 27628
rect 10100 27616 10106 27668
rect 10778 27616 10784 27668
rect 10836 27656 10842 27668
rect 11057 27659 11115 27665
rect 11057 27656 11069 27659
rect 10836 27628 11069 27656
rect 10836 27616 10842 27628
rect 11057 27625 11069 27628
rect 11103 27625 11115 27659
rect 11057 27619 11115 27625
rect 14182 27616 14188 27668
rect 14240 27616 14246 27668
rect 14734 27616 14740 27668
rect 14792 27656 14798 27668
rect 14829 27659 14887 27665
rect 14829 27656 14841 27659
rect 14792 27628 14841 27656
rect 14792 27616 14798 27628
rect 14829 27625 14841 27628
rect 14875 27625 14887 27659
rect 14829 27619 14887 27625
rect 15841 27659 15899 27665
rect 15841 27625 15853 27659
rect 15887 27656 15899 27659
rect 16114 27656 16120 27668
rect 15887 27628 16120 27656
rect 15887 27625 15899 27628
rect 15841 27619 15899 27625
rect 16114 27616 16120 27628
rect 16172 27616 16178 27668
rect 16390 27616 16396 27668
rect 16448 27656 16454 27668
rect 17862 27656 17868 27668
rect 16448 27628 17868 27656
rect 16448 27616 16454 27628
rect 17862 27616 17868 27628
rect 17920 27616 17926 27668
rect 18046 27616 18052 27668
rect 18104 27616 18110 27668
rect 18877 27659 18935 27665
rect 18877 27656 18889 27659
rect 18156 27628 18889 27656
rect 6362 27548 6368 27600
rect 6420 27588 6426 27600
rect 6546 27588 6552 27600
rect 6420 27560 6552 27588
rect 6420 27548 6426 27560
rect 6546 27548 6552 27560
rect 6604 27588 6610 27600
rect 6604 27560 7604 27588
rect 6604 27548 6610 27560
rect 3694 27480 3700 27532
rect 3752 27520 3758 27532
rect 4798 27520 4804 27532
rect 3752 27492 4804 27520
rect 3752 27480 3758 27492
rect 4798 27480 4804 27492
rect 4856 27480 4862 27532
rect 842 27412 848 27464
rect 900 27452 906 27464
rect 1397 27455 1455 27461
rect 1397 27452 1409 27455
rect 900 27424 1409 27452
rect 900 27412 906 27424
rect 1397 27421 1409 27424
rect 1443 27421 1455 27455
rect 1397 27415 1455 27421
rect 1670 27412 1676 27464
rect 1728 27412 1734 27464
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 6822 27452 6828 27464
rect 6512 27424 6828 27452
rect 6512 27412 6518 27424
rect 6822 27412 6828 27424
rect 6880 27452 6886 27464
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 6880 27424 7205 27452
rect 6880 27412 6886 27424
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 7193 27415 7251 27421
rect 7374 27412 7380 27464
rect 7432 27412 7438 27464
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 7576 27452 7604 27560
rect 10686 27548 10692 27600
rect 10744 27548 10750 27600
rect 13170 27548 13176 27600
rect 13228 27548 13234 27600
rect 17037 27591 17095 27597
rect 17037 27557 17049 27591
rect 17083 27588 17095 27591
rect 17126 27588 17132 27600
rect 17083 27560 17132 27588
rect 17083 27557 17095 27560
rect 17037 27551 17095 27557
rect 17126 27548 17132 27560
rect 17184 27548 17190 27600
rect 17497 27591 17555 27597
rect 17497 27557 17509 27591
rect 17543 27588 17555 27591
rect 17586 27588 17592 27600
rect 17543 27560 17592 27588
rect 17543 27557 17555 27560
rect 17497 27551 17555 27557
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 17770 27548 17776 27600
rect 17828 27588 17834 27600
rect 18156 27588 18184 27628
rect 18877 27625 18889 27628
rect 18923 27656 18935 27659
rect 18966 27656 18972 27668
rect 18923 27628 18972 27656
rect 18923 27625 18935 27628
rect 18877 27619 18935 27625
rect 18966 27616 18972 27628
rect 19024 27616 19030 27668
rect 19426 27616 19432 27668
rect 19484 27656 19490 27668
rect 19889 27659 19947 27665
rect 19889 27656 19901 27659
rect 19484 27628 19901 27656
rect 19484 27616 19490 27628
rect 19889 27625 19901 27628
rect 19935 27625 19947 27659
rect 19889 27619 19947 27625
rect 23587 27659 23645 27665
rect 23587 27625 23599 27659
rect 23633 27656 23645 27659
rect 23842 27656 23848 27668
rect 23633 27628 23848 27656
rect 23633 27625 23645 27628
rect 23587 27619 23645 27625
rect 23842 27616 23848 27628
rect 23900 27616 23906 27668
rect 25038 27616 25044 27668
rect 25096 27656 25102 27668
rect 25317 27659 25375 27665
rect 25317 27656 25329 27659
rect 25096 27628 25329 27656
rect 25096 27616 25102 27628
rect 25317 27625 25329 27628
rect 25363 27625 25375 27659
rect 25317 27619 25375 27625
rect 25774 27616 25780 27668
rect 25832 27616 25838 27668
rect 17828 27560 18184 27588
rect 19061 27591 19119 27597
rect 17828 27548 17834 27560
rect 19061 27557 19073 27591
rect 19107 27588 19119 27591
rect 19521 27591 19579 27597
rect 19521 27588 19533 27591
rect 19107 27560 19533 27588
rect 19107 27557 19119 27560
rect 19061 27551 19119 27557
rect 19521 27557 19533 27560
rect 19567 27588 19579 27591
rect 19610 27588 19616 27600
rect 19567 27560 19616 27588
rect 19567 27557 19579 27560
rect 19521 27551 19579 27557
rect 19610 27548 19616 27560
rect 19668 27548 19674 27600
rect 8021 27523 8079 27529
rect 8021 27489 8033 27523
rect 8067 27520 8079 27523
rect 8202 27520 8208 27532
rect 8067 27492 8208 27520
rect 8067 27489 8079 27492
rect 8021 27483 8079 27489
rect 8202 27480 8208 27492
rect 8260 27520 8266 27532
rect 10134 27520 10140 27532
rect 8260 27492 10140 27520
rect 8260 27480 8266 27492
rect 7745 27455 7803 27461
rect 7745 27452 7757 27455
rect 7576 27424 7757 27452
rect 7745 27421 7757 27424
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 8478 27412 8484 27464
rect 8536 27452 8542 27464
rect 8665 27455 8723 27461
rect 8665 27452 8677 27455
rect 8536 27424 8677 27452
rect 8536 27412 8542 27424
rect 8665 27421 8677 27424
rect 8711 27421 8723 27455
rect 8665 27415 8723 27421
rect 9122 27412 9128 27464
rect 9180 27412 9186 27464
rect 9876 27461 9904 27492
rect 10134 27480 10140 27492
rect 10192 27520 10198 27532
rect 10192 27492 13584 27520
rect 10192 27480 10198 27492
rect 9861 27455 9919 27461
rect 9861 27421 9873 27455
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 10042 27412 10048 27464
rect 10100 27452 10106 27464
rect 10226 27452 10232 27464
rect 10100 27424 10232 27452
rect 10100 27412 10106 27424
rect 10226 27412 10232 27424
rect 10284 27412 10290 27464
rect 11330 27412 11336 27464
rect 11388 27412 11394 27464
rect 13556 27461 13584 27492
rect 15010 27480 15016 27532
rect 15068 27520 15074 27532
rect 15068 27492 15516 27520
rect 15068 27480 15074 27492
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27421 13599 27455
rect 13541 27415 13599 27421
rect 13998 27412 14004 27464
rect 14056 27452 14062 27464
rect 14185 27455 14243 27461
rect 14185 27452 14197 27455
rect 14056 27424 14197 27452
rect 14056 27412 14062 27424
rect 14185 27421 14197 27424
rect 14231 27421 14243 27455
rect 14185 27415 14243 27421
rect 14366 27412 14372 27464
rect 14424 27412 14430 27464
rect 14461 27455 14519 27461
rect 14461 27421 14473 27455
rect 14507 27452 14519 27455
rect 14826 27452 14832 27464
rect 14507 27424 14832 27452
rect 14507 27421 14519 27424
rect 14461 27415 14519 27421
rect 5077 27387 5135 27393
rect 5077 27353 5089 27387
rect 5123 27384 5135 27387
rect 5350 27384 5356 27396
rect 5123 27356 5356 27384
rect 5123 27353 5135 27356
rect 5077 27347 5135 27353
rect 5350 27344 5356 27356
rect 5408 27344 5414 27396
rect 5810 27344 5816 27396
rect 5868 27344 5874 27396
rect 6362 27344 6368 27396
rect 6420 27384 6426 27396
rect 6917 27387 6975 27393
rect 6917 27384 6929 27387
rect 6420 27356 6929 27384
rect 6420 27344 6426 27356
rect 6917 27353 6929 27356
rect 6963 27353 6975 27387
rect 6917 27347 6975 27353
rect 7098 27344 7104 27396
rect 7156 27344 7162 27396
rect 7834 27344 7840 27396
rect 7892 27344 7898 27396
rect 8018 27344 8024 27396
rect 8076 27384 8082 27396
rect 8297 27387 8355 27393
rect 8297 27384 8309 27387
rect 8076 27356 8309 27384
rect 8076 27344 8082 27356
rect 8297 27353 8309 27356
rect 8343 27353 8355 27387
rect 9140 27384 9168 27412
rect 10962 27384 10968 27396
rect 9140 27356 10968 27384
rect 8297 27347 8355 27353
rect 10962 27344 10968 27356
rect 11020 27344 11026 27396
rect 11054 27344 11060 27396
rect 11112 27344 11118 27396
rect 11609 27387 11667 27393
rect 11609 27353 11621 27387
rect 11655 27353 11667 27387
rect 11609 27347 11667 27353
rect 6638 27276 6644 27328
rect 6696 27316 6702 27328
rect 6733 27319 6791 27325
rect 6733 27316 6745 27319
rect 6696 27288 6745 27316
rect 6696 27276 6702 27288
rect 6733 27285 6745 27288
rect 6779 27285 6791 27319
rect 6733 27279 6791 27285
rect 7650 27276 7656 27328
rect 7708 27276 7714 27328
rect 8110 27276 8116 27328
rect 8168 27276 8174 27328
rect 9033 27319 9091 27325
rect 9033 27285 9045 27319
rect 9079 27316 9091 27319
rect 9122 27316 9128 27328
rect 9079 27288 9128 27316
rect 9079 27285 9091 27288
rect 9033 27279 9091 27285
rect 9122 27276 9128 27288
rect 9180 27276 9186 27328
rect 11241 27319 11299 27325
rect 11241 27285 11253 27319
rect 11287 27316 11299 27319
rect 11624 27316 11652 27347
rect 12618 27344 12624 27396
rect 12676 27344 12682 27396
rect 13725 27387 13783 27393
rect 13725 27353 13737 27387
rect 13771 27384 13783 27387
rect 14090 27384 14096 27396
rect 13771 27356 14096 27384
rect 13771 27353 13783 27356
rect 13725 27347 13783 27353
rect 14090 27344 14096 27356
rect 14148 27384 14154 27396
rect 14476 27384 14504 27415
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 15105 27455 15163 27461
rect 15105 27421 15117 27455
rect 15151 27452 15163 27455
rect 15378 27452 15384 27464
rect 15151 27424 15384 27452
rect 15151 27421 15163 27424
rect 15105 27415 15163 27421
rect 14148 27356 14504 27384
rect 14645 27387 14703 27393
rect 14148 27344 14154 27356
rect 14645 27353 14657 27387
rect 14691 27384 14703 27387
rect 15120 27384 15148 27415
rect 15378 27412 15384 27424
rect 15436 27412 15442 27464
rect 15488 27461 15516 27492
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27421 15531 27455
rect 15473 27415 15531 27421
rect 16942 27412 16948 27464
rect 17000 27412 17006 27464
rect 17604 27452 17632 27548
rect 19978 27480 19984 27532
rect 20036 27520 20042 27532
rect 20165 27523 20223 27529
rect 20165 27520 20177 27523
rect 20036 27492 20177 27520
rect 20036 27480 20042 27492
rect 20165 27489 20177 27492
rect 20211 27489 20223 27523
rect 20165 27483 20223 27489
rect 22097 27523 22155 27529
rect 22097 27489 22109 27523
rect 22143 27520 22155 27523
rect 23474 27520 23480 27532
rect 22143 27492 23480 27520
rect 22143 27489 22155 27492
rect 22097 27483 22155 27489
rect 23474 27480 23480 27492
rect 23532 27480 23538 27532
rect 17604 27424 18828 27452
rect 14691 27356 15148 27384
rect 14691 27353 14703 27356
rect 14645 27347 14703 27353
rect 15286 27344 15292 27396
rect 15344 27384 15350 27396
rect 15562 27384 15568 27396
rect 15344 27356 15568 27384
rect 15344 27344 15350 27356
rect 15562 27344 15568 27356
rect 15620 27384 15626 27396
rect 15657 27387 15715 27393
rect 15657 27384 15669 27387
rect 15620 27356 15669 27384
rect 15620 27344 15626 27356
rect 15657 27353 15669 27356
rect 15703 27384 15715 27387
rect 16758 27384 16764 27396
rect 15703 27356 16764 27384
rect 15703 27353 15715 27356
rect 15657 27347 15715 27353
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 17865 27387 17923 27393
rect 17865 27353 17877 27387
rect 17911 27384 17923 27387
rect 17954 27384 17960 27396
rect 17911 27356 17960 27384
rect 17911 27353 17923 27356
rect 17865 27347 17923 27353
rect 17954 27344 17960 27356
rect 18012 27344 18018 27396
rect 18693 27387 18751 27393
rect 18693 27353 18705 27387
rect 18739 27353 18751 27387
rect 18800 27384 18828 27424
rect 19242 27412 19248 27464
rect 19300 27412 19306 27464
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27452 19487 27455
rect 19702 27452 19708 27464
rect 19475 27424 19708 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 19702 27412 19708 27424
rect 19760 27412 19766 27464
rect 23845 27455 23903 27461
rect 23845 27421 23857 27455
rect 23891 27452 23903 27455
rect 24762 27452 24768 27464
rect 23891 27424 24768 27452
rect 23891 27421 23903 27424
rect 23845 27415 23903 27421
rect 24762 27412 24768 27424
rect 24820 27412 24826 27464
rect 25130 27412 25136 27464
rect 25188 27412 25194 27464
rect 25314 27412 25320 27464
rect 25372 27412 25378 27464
rect 27062 27412 27068 27464
rect 27120 27452 27126 27464
rect 27614 27452 27620 27464
rect 27120 27424 27620 27452
rect 27120 27412 27126 27424
rect 27614 27412 27620 27424
rect 27672 27412 27678 27464
rect 18893 27387 18951 27393
rect 18893 27384 18905 27387
rect 18800 27356 18905 27384
rect 18693 27347 18751 27353
rect 18893 27353 18905 27356
rect 18939 27353 18951 27387
rect 20441 27387 20499 27393
rect 20441 27384 20453 27387
rect 18893 27347 18951 27353
rect 20088 27356 20453 27384
rect 11287 27288 11652 27316
rect 13081 27319 13139 27325
rect 11287 27285 11299 27288
rect 11241 27279 11299 27285
rect 13081 27285 13093 27319
rect 13127 27316 13139 27319
rect 13262 27316 13268 27328
rect 13127 27288 13268 27316
rect 13127 27285 13139 27288
rect 13081 27279 13139 27285
rect 13262 27276 13268 27288
rect 13320 27316 13326 27328
rect 13357 27319 13415 27325
rect 13357 27316 13369 27319
rect 13320 27288 13369 27316
rect 13320 27276 13326 27288
rect 13357 27285 13369 27288
rect 13403 27285 13415 27319
rect 13357 27279 13415 27285
rect 13449 27319 13507 27325
rect 13449 27285 13461 27319
rect 13495 27316 13507 27319
rect 13538 27316 13544 27328
rect 13495 27288 13544 27316
rect 13495 27285 13507 27288
rect 13449 27279 13507 27285
rect 13538 27276 13544 27288
rect 13596 27276 13602 27328
rect 14182 27276 14188 27328
rect 14240 27316 14246 27328
rect 14366 27316 14372 27328
rect 14240 27288 14372 27316
rect 14240 27276 14246 27288
rect 14366 27276 14372 27288
rect 14424 27316 14430 27328
rect 15013 27319 15071 27325
rect 15013 27316 15025 27319
rect 14424 27288 15025 27316
rect 14424 27276 14430 27288
rect 15013 27285 15025 27288
rect 15059 27285 15071 27319
rect 18708 27316 18736 27347
rect 19334 27316 19340 27328
rect 18708 27288 19340 27316
rect 15013 27279 15071 27285
rect 19334 27276 19340 27288
rect 19392 27276 19398 27328
rect 20088 27325 20116 27356
rect 20441 27353 20453 27356
rect 20487 27353 20499 27387
rect 20441 27347 20499 27353
rect 21174 27344 21180 27396
rect 21232 27344 21238 27396
rect 22554 27344 22560 27396
rect 22612 27344 22618 27396
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 19889 27319 19947 27325
rect 19889 27316 19901 27319
rect 19475 27288 19901 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 19889 27285 19901 27288
rect 19935 27285 19947 27319
rect 19889 27279 19947 27285
rect 20073 27319 20131 27325
rect 20073 27285 20085 27319
rect 20119 27285 20131 27319
rect 20073 27279 20131 27285
rect 20622 27276 20628 27328
rect 20680 27316 20686 27328
rect 21913 27319 21971 27325
rect 21913 27316 21925 27319
rect 20680 27288 21925 27316
rect 20680 27276 20686 27288
rect 21913 27285 21925 27288
rect 21959 27285 21971 27319
rect 25148 27316 25176 27412
rect 25498 27344 25504 27396
rect 25556 27384 25562 27396
rect 25745 27387 25803 27393
rect 25745 27384 25757 27387
rect 25556 27356 25757 27384
rect 25556 27344 25562 27356
rect 25745 27353 25757 27356
rect 25791 27384 25803 27387
rect 25866 27384 25872 27396
rect 25791 27356 25872 27384
rect 25791 27353 25803 27356
rect 25745 27347 25803 27353
rect 25866 27344 25872 27356
rect 25924 27344 25930 27396
rect 25958 27344 25964 27396
rect 26016 27344 26022 27396
rect 27890 27344 27896 27396
rect 27948 27344 27954 27396
rect 28902 27344 28908 27396
rect 28960 27344 28966 27396
rect 25593 27319 25651 27325
rect 25593 27316 25605 27319
rect 25148 27288 25605 27316
rect 21913 27279 21971 27285
rect 25593 27285 25605 27288
rect 25639 27285 25651 27319
rect 25593 27279 25651 27285
rect 27982 27276 27988 27328
rect 28040 27316 28046 27328
rect 29365 27319 29423 27325
rect 29365 27316 29377 27319
rect 28040 27288 29377 27316
rect 28040 27276 28046 27288
rect 29365 27285 29377 27288
rect 29411 27285 29423 27319
rect 29365 27279 29423 27285
rect 1104 27226 29716 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 29716 27226
rect 1104 27152 29716 27174
rect 5350 27072 5356 27124
rect 5408 27112 5414 27124
rect 6365 27115 6423 27121
rect 6365 27112 6377 27115
rect 5408 27084 6377 27112
rect 5408 27072 5414 27084
rect 6365 27081 6377 27084
rect 6411 27081 6423 27115
rect 6365 27075 6423 27081
rect 6533 27115 6591 27121
rect 6533 27081 6545 27115
rect 6579 27112 6591 27115
rect 6638 27112 6644 27124
rect 6579 27084 6644 27112
rect 6579 27081 6591 27084
rect 6533 27075 6591 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7009 27115 7067 27121
rect 7009 27081 7021 27115
rect 7055 27112 7067 27115
rect 7558 27112 7564 27124
rect 7055 27084 7564 27112
rect 7055 27081 7067 27084
rect 7009 27075 7067 27081
rect 7558 27072 7564 27084
rect 7616 27112 7622 27124
rect 8478 27112 8484 27124
rect 7616 27084 8484 27112
rect 7616 27072 7622 27084
rect 8478 27072 8484 27084
rect 8536 27072 8542 27124
rect 9582 27072 9588 27124
rect 9640 27072 9646 27124
rect 12437 27115 12495 27121
rect 12437 27081 12449 27115
rect 12483 27112 12495 27115
rect 12618 27112 12624 27124
rect 12483 27084 12624 27112
rect 12483 27081 12495 27084
rect 12437 27075 12495 27081
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 13998 27072 14004 27124
rect 14056 27072 14062 27124
rect 18506 27072 18512 27124
rect 18564 27072 18570 27124
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 20622 27112 20628 27124
rect 19392 27084 20628 27112
rect 19392 27072 19398 27084
rect 20622 27072 20628 27084
rect 20680 27072 20686 27124
rect 21174 27072 21180 27124
rect 21232 27112 21238 27124
rect 21269 27115 21327 27121
rect 21269 27112 21281 27115
rect 21232 27084 21281 27112
rect 21232 27072 21238 27084
rect 21269 27081 21281 27084
rect 21315 27081 21327 27115
rect 21269 27075 21327 27081
rect 22554 27072 22560 27124
rect 22612 27112 22618 27124
rect 22649 27115 22707 27121
rect 22649 27112 22661 27115
rect 22612 27084 22661 27112
rect 22612 27072 22618 27084
rect 22649 27081 22661 27084
rect 22695 27081 22707 27115
rect 22649 27075 22707 27081
rect 27709 27115 27767 27121
rect 27709 27081 27721 27115
rect 27755 27112 27767 27115
rect 27890 27112 27896 27124
rect 27755 27084 27896 27112
rect 27755 27081 27767 27084
rect 27709 27075 27767 27081
rect 27890 27072 27896 27084
rect 27948 27072 27954 27124
rect 28902 27072 28908 27124
rect 28960 27072 28966 27124
rect 6178 27004 6184 27056
rect 6236 27044 6242 27056
rect 6733 27047 6791 27053
rect 6733 27044 6745 27047
rect 6236 27016 6745 27044
rect 6236 27004 6242 27016
rect 6733 27013 6745 27016
rect 6779 27013 6791 27047
rect 6733 27007 6791 27013
rect 6748 26908 6776 27007
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 6880 27016 7144 27044
rect 6880 27004 6886 27016
rect 6914 26936 6920 26988
rect 6972 26936 6978 26988
rect 7116 26985 7144 27016
rect 7282 27004 7288 27056
rect 7340 27044 7346 27056
rect 8018 27044 8024 27056
rect 7340 27016 8024 27044
rect 7340 27004 7346 27016
rect 8018 27004 8024 27016
rect 8076 27004 8082 27056
rect 8110 27004 8116 27056
rect 8168 27004 8174 27056
rect 9122 27004 9128 27056
rect 9180 27004 9186 27056
rect 9600 27044 9628 27072
rect 18524 27044 18552 27072
rect 19242 27044 19248 27056
rect 9600 27016 9674 27044
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26945 7159 26979
rect 7101 26939 7159 26945
rect 7300 26908 7328 27004
rect 7742 26936 7748 26988
rect 7800 26976 7806 26988
rect 7837 26979 7895 26985
rect 7837 26976 7849 26979
rect 7800 26948 7849 26976
rect 7800 26936 7806 26948
rect 7837 26945 7849 26948
rect 7883 26945 7895 26979
rect 9646 26976 9674 27016
rect 10428 27016 19248 27044
rect 9769 26979 9827 26985
rect 9769 26976 9781 26979
rect 9646 26948 9781 26976
rect 7837 26939 7895 26945
rect 9769 26945 9781 26948
rect 9815 26945 9827 26979
rect 9769 26939 9827 26945
rect 6748 26880 7328 26908
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 9861 26911 9919 26917
rect 9861 26908 9873 26911
rect 7432 26880 9873 26908
rect 7432 26868 7438 26880
rect 9861 26877 9873 26880
rect 9907 26908 9919 26911
rect 10318 26908 10324 26920
rect 9907 26880 10324 26908
rect 9907 26877 9919 26880
rect 9861 26871 9919 26877
rect 10318 26868 10324 26880
rect 10376 26868 10382 26920
rect 3326 26800 3332 26852
rect 3384 26840 3390 26852
rect 10428 26840 10456 27016
rect 19242 27004 19248 27016
rect 19300 27004 19306 27056
rect 24486 27004 24492 27056
rect 24544 27004 24550 27056
rect 29270 27004 29276 27056
rect 29328 27004 29334 27056
rect 10962 26936 10968 26988
rect 11020 26976 11026 26988
rect 12345 26979 12403 26985
rect 12345 26976 12357 26979
rect 11020 26948 12357 26976
rect 11020 26936 11026 26948
rect 12345 26945 12357 26948
rect 12391 26976 12403 26979
rect 12434 26976 12440 26988
rect 12391 26948 12440 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 13262 26936 13268 26988
rect 13320 26936 13326 26988
rect 14090 26936 14096 26988
rect 14148 26936 14154 26988
rect 14826 26936 14832 26988
rect 14884 26936 14890 26988
rect 15197 26979 15255 26985
rect 15197 26945 15209 26979
rect 15243 26976 15255 26979
rect 15930 26976 15936 26988
rect 15243 26948 15936 26976
rect 15243 26945 15255 26948
rect 15197 26939 15255 26945
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 18509 26979 18567 26985
rect 18509 26945 18521 26979
rect 18555 26976 18567 26979
rect 18598 26976 18604 26988
rect 18555 26948 18604 26976
rect 18555 26945 18567 26948
rect 18509 26939 18567 26945
rect 18598 26936 18604 26948
rect 18656 26936 18662 26988
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 21082 26936 21088 26988
rect 21140 26976 21146 26988
rect 21177 26979 21235 26985
rect 21177 26976 21189 26979
rect 21140 26948 21189 26976
rect 21140 26936 21146 26948
rect 21177 26945 21189 26948
rect 21223 26976 21235 26979
rect 22002 26976 22008 26988
rect 21223 26948 22008 26976
rect 21223 26945 21235 26948
rect 21177 26939 21235 26945
rect 22002 26936 22008 26948
rect 22060 26976 22066 26988
rect 22557 26979 22615 26985
rect 22557 26976 22569 26979
rect 22060 26948 22569 26976
rect 22060 26936 22066 26948
rect 22557 26945 22569 26948
rect 22603 26945 22615 26979
rect 22557 26939 22615 26945
rect 25225 26979 25283 26985
rect 25225 26945 25237 26979
rect 25271 26976 25283 26979
rect 27062 26976 27068 26988
rect 25271 26948 27068 26976
rect 25271 26945 25283 26948
rect 25225 26939 25283 26945
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 13357 26911 13415 26917
rect 13357 26908 13369 26911
rect 11204 26880 13369 26908
rect 11204 26868 11210 26880
rect 13357 26877 13369 26880
rect 13403 26908 13415 26911
rect 13722 26908 13728 26920
rect 13403 26880 13728 26908
rect 13403 26877 13415 26880
rect 13357 26871 13415 26877
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 23474 26868 23480 26920
rect 23532 26908 23538 26920
rect 23750 26908 23756 26920
rect 23532 26880 23756 26908
rect 23532 26868 23538 26880
rect 23750 26868 23756 26880
rect 23808 26868 23814 26920
rect 24946 26868 24952 26920
rect 25004 26868 25010 26920
rect 3384 26812 7972 26840
rect 3384 26800 3390 26812
rect 6549 26775 6607 26781
rect 6549 26741 6561 26775
rect 6595 26772 6607 26775
rect 6822 26772 6828 26784
rect 6595 26744 6828 26772
rect 6595 26741 6607 26744
rect 6549 26735 6607 26741
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 6914 26732 6920 26784
rect 6972 26772 6978 26784
rect 7374 26772 7380 26784
rect 6972 26744 7380 26772
rect 6972 26732 6978 26744
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 7944 26772 7972 26812
rect 9508 26812 10456 26840
rect 9508 26772 9536 26812
rect 12618 26800 12624 26852
rect 12676 26840 12682 26852
rect 13446 26840 13452 26852
rect 12676 26812 13452 26840
rect 12676 26800 12682 26812
rect 13446 26800 13452 26812
rect 13504 26800 13510 26852
rect 17862 26800 17868 26852
rect 17920 26840 17926 26852
rect 18414 26840 18420 26852
rect 17920 26812 18420 26840
rect 17920 26800 17926 26812
rect 18414 26800 18420 26812
rect 18472 26840 18478 26852
rect 20714 26840 20720 26852
rect 18472 26812 20720 26840
rect 18472 26800 18478 26812
rect 20714 26800 20720 26812
rect 20772 26800 20778 26852
rect 7944 26744 9536 26772
rect 10042 26732 10048 26784
rect 10100 26772 10106 26784
rect 13170 26772 13176 26784
rect 10100 26744 13176 26772
rect 10100 26732 10106 26744
rect 13170 26732 13176 26744
rect 13228 26772 13234 26784
rect 13538 26772 13544 26784
rect 13228 26744 13544 26772
rect 13228 26732 13234 26744
rect 13538 26732 13544 26744
rect 13596 26732 13602 26784
rect 15194 26732 15200 26784
rect 15252 26732 15258 26784
rect 15286 26732 15292 26784
rect 15344 26772 15350 26784
rect 15381 26775 15439 26781
rect 15381 26772 15393 26775
rect 15344 26744 15393 26772
rect 15344 26732 15350 26744
rect 15381 26741 15393 26744
rect 15427 26741 15439 26775
rect 15381 26735 15439 26741
rect 15746 26732 15752 26784
rect 15804 26772 15810 26784
rect 18509 26775 18567 26781
rect 18509 26772 18521 26775
rect 15804 26744 18521 26772
rect 15804 26732 15810 26744
rect 18509 26741 18521 26744
rect 18555 26741 18567 26775
rect 18509 26735 18567 26741
rect 23474 26732 23480 26784
rect 23532 26732 23538 26784
rect 24762 26732 24768 26784
rect 24820 26772 24826 26784
rect 25240 26772 25268 26939
rect 27062 26936 27068 26948
rect 27120 26936 27126 26988
rect 27341 26979 27399 26985
rect 27341 26945 27353 26979
rect 27387 26976 27399 26979
rect 27982 26976 27988 26988
rect 27387 26948 27988 26976
rect 27387 26945 27399 26948
rect 27341 26939 27399 26945
rect 27982 26936 27988 26948
rect 28040 26936 28046 26988
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26976 29055 26979
rect 29086 26976 29092 26988
rect 29043 26948 29092 26976
rect 29043 26945 29055 26948
rect 28997 26939 29055 26945
rect 29086 26936 29092 26948
rect 29144 26936 29150 26988
rect 27430 26868 27436 26920
rect 27488 26868 27494 26920
rect 24820 26744 25268 26772
rect 29181 26775 29239 26781
rect 24820 26732 24826 26744
rect 29181 26741 29193 26775
rect 29227 26772 29239 26775
rect 29546 26772 29552 26784
rect 29227 26744 29552 26772
rect 29227 26741 29239 26744
rect 29181 26735 29239 26741
rect 29546 26732 29552 26744
rect 29604 26732 29610 26784
rect 1104 26682 29716 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 29716 26682
rect 1104 26608 29716 26630
rect 16850 26568 16856 26580
rect 6472 26540 16856 26568
rect 4798 26432 4804 26444
rect 4264 26404 4804 26432
rect 4264 26373 4292 26404
rect 4798 26392 4804 26404
rect 4856 26392 4862 26444
rect 4249 26367 4307 26373
rect 4249 26333 4261 26367
rect 4295 26333 4307 26367
rect 4706 26364 4712 26376
rect 4249 26327 4307 26333
rect 4356 26336 4712 26364
rect 1486 26256 1492 26308
rect 1544 26256 1550 26308
rect 1673 26299 1731 26305
rect 1673 26265 1685 26299
rect 1719 26296 1731 26299
rect 2038 26296 2044 26308
rect 1719 26268 2044 26296
rect 1719 26265 1731 26268
rect 1673 26259 1731 26265
rect 2038 26256 2044 26268
rect 2096 26256 2102 26308
rect 4154 26256 4160 26308
rect 4212 26296 4218 26308
rect 4356 26296 4384 26336
rect 4706 26324 4712 26336
rect 4764 26324 4770 26376
rect 6472 26373 6500 26540
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 18049 26571 18107 26577
rect 18049 26568 18061 26571
rect 16960 26540 18061 26568
rect 11149 26503 11207 26509
rect 11149 26469 11161 26503
rect 11195 26500 11207 26503
rect 12618 26500 12624 26512
rect 11195 26472 12624 26500
rect 11195 26469 11207 26472
rect 11149 26463 11207 26469
rect 12618 26460 12624 26472
rect 12676 26460 12682 26512
rect 16025 26503 16083 26509
rect 12728 26472 13400 26500
rect 8478 26392 8484 26444
rect 8536 26432 8542 26444
rect 8536 26404 11652 26432
rect 8536 26392 8542 26404
rect 6457 26367 6515 26373
rect 5184 26336 6408 26364
rect 4212 26268 4384 26296
rect 4433 26299 4491 26305
rect 4212 26256 4218 26268
rect 4433 26265 4445 26299
rect 4479 26296 4491 26299
rect 5184 26296 5212 26336
rect 4479 26268 5212 26296
rect 4479 26265 4491 26268
rect 4433 26259 4491 26265
rect 4614 26188 4620 26240
rect 4672 26188 4678 26240
rect 4706 26188 4712 26240
rect 4764 26228 4770 26240
rect 4801 26231 4859 26237
rect 4801 26228 4813 26231
rect 4764 26200 4813 26228
rect 4764 26188 4770 26200
rect 4801 26197 4813 26200
rect 4847 26197 4859 26231
rect 5184 26228 5212 26268
rect 5258 26256 5264 26308
rect 5316 26296 5322 26308
rect 5813 26299 5871 26305
rect 5813 26296 5825 26299
rect 5316 26268 5825 26296
rect 5316 26256 5322 26268
rect 5813 26265 5825 26268
rect 5859 26265 5871 26299
rect 5813 26259 5871 26265
rect 5994 26256 6000 26308
rect 6052 26256 6058 26308
rect 6380 26296 6408 26336
rect 6457 26333 6469 26367
rect 6503 26364 6515 26367
rect 6638 26364 6644 26376
rect 6503 26336 6644 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 6638 26324 6644 26336
rect 6696 26324 6702 26376
rect 6733 26367 6791 26373
rect 6733 26333 6745 26367
rect 6779 26333 6791 26367
rect 6733 26327 6791 26333
rect 8389 26367 8447 26373
rect 8389 26333 8401 26367
rect 8435 26364 8447 26367
rect 8570 26364 8576 26376
rect 8435 26336 8576 26364
rect 8435 26333 8447 26336
rect 8389 26327 8447 26333
rect 6748 26296 6776 26327
rect 8570 26324 8576 26336
rect 8628 26324 8634 26376
rect 9398 26324 9404 26376
rect 9456 26324 9462 26376
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9508 26296 9536 26327
rect 10134 26324 10140 26376
rect 10192 26324 10198 26376
rect 10318 26324 10324 26376
rect 10376 26324 10382 26376
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26364 10563 26367
rect 11238 26364 11244 26376
rect 10551 26336 11244 26364
rect 10551 26333 10563 26336
rect 10505 26327 10563 26333
rect 11238 26324 11244 26336
rect 11296 26364 11302 26376
rect 11333 26367 11391 26373
rect 11333 26364 11345 26367
rect 11296 26336 11345 26364
rect 11296 26324 11302 26336
rect 11333 26333 11345 26336
rect 11379 26333 11391 26367
rect 11333 26327 11391 26333
rect 11425 26367 11483 26373
rect 11425 26333 11437 26367
rect 11471 26333 11483 26367
rect 11425 26327 11483 26333
rect 11624 26364 11652 26404
rect 11698 26392 11704 26444
rect 11756 26432 11762 26444
rect 11793 26435 11851 26441
rect 11793 26432 11805 26435
rect 11756 26404 11805 26432
rect 11756 26392 11762 26404
rect 11793 26401 11805 26404
rect 11839 26432 11851 26435
rect 12728 26432 12756 26472
rect 11839 26404 12756 26432
rect 11839 26401 11851 26404
rect 11793 26395 11851 26401
rect 12728 26373 12756 26404
rect 13170 26392 13176 26444
rect 13228 26392 13234 26444
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 11624 26336 12633 26364
rect 6380 26268 6776 26296
rect 8312 26268 9536 26296
rect 10152 26296 10180 26324
rect 10152 26268 10548 26296
rect 8312 26240 8340 26268
rect 5350 26228 5356 26240
rect 5184 26200 5356 26228
rect 4801 26191 4859 26197
rect 5350 26188 5356 26200
rect 5408 26188 5414 26240
rect 6181 26231 6239 26237
rect 6181 26197 6193 26231
rect 6227 26228 6239 26231
rect 6270 26228 6276 26240
rect 6227 26200 6276 26228
rect 6227 26197 6239 26200
rect 6181 26191 6239 26197
rect 6270 26188 6276 26200
rect 6328 26188 6334 26240
rect 6365 26231 6423 26237
rect 6365 26197 6377 26231
rect 6411 26228 6423 26231
rect 6454 26228 6460 26240
rect 6411 26200 6460 26228
rect 6411 26197 6423 26200
rect 6365 26191 6423 26197
rect 6454 26188 6460 26200
rect 6512 26188 6518 26240
rect 6641 26231 6699 26237
rect 6641 26197 6653 26231
rect 6687 26228 6699 26231
rect 6730 26228 6736 26240
rect 6687 26200 6736 26228
rect 6687 26197 6699 26200
rect 6641 26191 6699 26197
rect 6730 26188 6736 26200
rect 6788 26188 6794 26240
rect 7190 26188 7196 26240
rect 7248 26228 7254 26240
rect 7650 26228 7656 26240
rect 7248 26200 7656 26228
rect 7248 26188 7254 26200
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 8294 26188 8300 26240
rect 8352 26188 8358 26240
rect 9677 26231 9735 26237
rect 9677 26197 9689 26231
rect 9723 26228 9735 26231
rect 9858 26228 9864 26240
rect 9723 26200 9864 26228
rect 9723 26197 9735 26200
rect 9677 26191 9735 26197
rect 9858 26188 9864 26200
rect 9916 26188 9922 26240
rect 10520 26228 10548 26268
rect 10594 26256 10600 26308
rect 10652 26256 10658 26308
rect 10781 26299 10839 26305
rect 10781 26296 10793 26299
rect 10704 26268 10793 26296
rect 10704 26228 10732 26268
rect 10781 26265 10793 26268
rect 10827 26265 10839 26299
rect 10781 26259 10839 26265
rect 10870 26256 10876 26308
rect 10928 26296 10934 26308
rect 11440 26296 11468 26327
rect 10928 26268 11468 26296
rect 11624 26296 11652 26336
rect 12621 26333 12633 26336
rect 12667 26333 12679 26367
rect 12621 26327 12679 26333
rect 12713 26367 12771 26373
rect 12713 26333 12725 26367
rect 12759 26333 12771 26367
rect 12713 26327 12771 26333
rect 11701 26299 11759 26305
rect 11701 26296 11713 26299
rect 11624 26268 11713 26296
rect 10928 26256 10934 26268
rect 11701 26265 11713 26268
rect 11747 26265 11759 26299
rect 12636 26296 12664 26327
rect 12894 26324 12900 26376
rect 12952 26324 12958 26376
rect 12986 26324 12992 26376
rect 13044 26324 13050 26376
rect 13078 26324 13084 26376
rect 13136 26324 13142 26376
rect 13372 26373 13400 26472
rect 16025 26469 16037 26503
rect 16071 26469 16083 26503
rect 16025 26463 16083 26469
rect 14642 26392 14648 26444
rect 14700 26392 14706 26444
rect 13357 26367 13415 26373
rect 13357 26333 13369 26367
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 13449 26367 13507 26373
rect 13449 26333 13461 26367
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26333 15163 26367
rect 15105 26327 15163 26333
rect 13464 26296 13492 26327
rect 15120 26296 15148 26327
rect 15286 26324 15292 26376
rect 15344 26324 15350 26376
rect 15657 26367 15715 26373
rect 15657 26333 15669 26367
rect 15703 26364 15715 26367
rect 15746 26364 15752 26376
rect 15703 26336 15752 26364
rect 15703 26333 15715 26336
rect 15657 26327 15715 26333
rect 15746 26324 15752 26336
rect 15804 26324 15810 26376
rect 15841 26367 15899 26373
rect 15841 26333 15853 26367
rect 15887 26364 15899 26367
rect 16040 26364 16068 26463
rect 16960 26432 16988 26540
rect 18049 26537 18061 26540
rect 18095 26537 18107 26571
rect 18049 26531 18107 26537
rect 20257 26571 20315 26577
rect 20257 26537 20269 26571
rect 20303 26568 20315 26571
rect 20533 26571 20591 26577
rect 20533 26568 20545 26571
rect 20303 26540 20545 26568
rect 20303 26537 20315 26540
rect 20257 26531 20315 26537
rect 20533 26537 20545 26540
rect 20579 26537 20591 26571
rect 20533 26531 20591 26537
rect 20640 26540 23612 26568
rect 17126 26460 17132 26512
rect 17184 26500 17190 26512
rect 20640 26500 20668 26540
rect 17184 26472 20668 26500
rect 20717 26503 20775 26509
rect 17184 26460 17190 26472
rect 20717 26469 20729 26503
rect 20763 26500 20775 26503
rect 23290 26500 23296 26512
rect 20763 26472 23296 26500
rect 20763 26469 20775 26472
rect 20717 26463 20775 26469
rect 23290 26460 23296 26472
rect 23348 26460 23354 26512
rect 23477 26503 23535 26509
rect 23477 26469 23489 26503
rect 23523 26469 23535 26503
rect 23584 26500 23612 26540
rect 23750 26528 23756 26580
rect 23808 26528 23814 26580
rect 24029 26571 24087 26577
rect 24029 26537 24041 26571
rect 24075 26568 24087 26571
rect 24946 26568 24952 26580
rect 24075 26540 24952 26568
rect 24075 26537 24087 26540
rect 24029 26531 24087 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 29181 26571 29239 26577
rect 29181 26568 29193 26571
rect 25056 26540 29193 26568
rect 25056 26500 25084 26540
rect 29181 26537 29193 26540
rect 29227 26537 29239 26571
rect 29181 26531 29239 26537
rect 27433 26503 27491 26509
rect 27433 26500 27445 26503
rect 23584 26472 25084 26500
rect 26436 26472 27445 26500
rect 23477 26463 23535 26469
rect 16316 26404 16988 26432
rect 16316 26373 16344 26404
rect 17218 26392 17224 26444
rect 17276 26392 17282 26444
rect 18233 26435 18291 26441
rect 18233 26432 18245 26435
rect 17328 26404 18245 26432
rect 15887 26336 16068 26364
rect 16301 26367 16359 26373
rect 15887 26333 15899 26336
rect 15841 26327 15899 26333
rect 16301 26333 16313 26367
rect 16347 26333 16359 26367
rect 16301 26327 16359 26333
rect 16942 26324 16948 26376
rect 17000 26324 17006 26376
rect 17034 26324 17040 26376
rect 17092 26324 17098 26376
rect 17328 26373 17356 26404
rect 17512 26373 17540 26404
rect 18233 26401 18245 26404
rect 18279 26401 18291 26435
rect 19337 26435 19395 26441
rect 19337 26432 19349 26435
rect 18233 26395 18291 26401
rect 18708 26404 19349 26432
rect 18708 26376 18736 26404
rect 19337 26401 19349 26404
rect 19383 26401 19395 26435
rect 19337 26395 19395 26401
rect 19536 26404 19840 26432
rect 17313 26367 17371 26373
rect 17313 26333 17325 26367
rect 17359 26333 17371 26367
rect 17313 26327 17371 26333
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 17498 26367 17556 26373
rect 17498 26333 17510 26367
rect 17544 26364 17556 26367
rect 17911 26367 17969 26373
rect 17544 26336 17577 26364
rect 17544 26333 17556 26336
rect 17498 26327 17556 26333
rect 17911 26333 17923 26367
rect 17957 26364 17969 26367
rect 18046 26364 18052 26376
rect 17957 26336 18052 26364
rect 17957 26333 17969 26336
rect 17911 26327 17969 26333
rect 12636 26268 13492 26296
rect 13556 26268 15148 26296
rect 16025 26299 16083 26305
rect 11701 26259 11759 26265
rect 10520 26200 10732 26228
rect 10962 26188 10968 26240
rect 11020 26188 11026 26240
rect 12434 26188 12440 26240
rect 12492 26188 12498 26240
rect 12710 26188 12716 26240
rect 12768 26228 12774 26240
rect 13556 26228 13584 26268
rect 16025 26265 16037 26299
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 12768 26200 13584 26228
rect 12768 26188 12774 26200
rect 13630 26188 13636 26240
rect 13688 26188 13694 26240
rect 16040 26228 16068 26259
rect 16206 26256 16212 26308
rect 16264 26256 16270 26308
rect 16761 26299 16819 26305
rect 16761 26265 16773 26299
rect 16807 26296 16819 26299
rect 17420 26296 17448 26327
rect 18046 26324 18052 26336
rect 18104 26364 18110 26376
rect 18325 26367 18383 26373
rect 18104 26336 18276 26364
rect 18104 26324 18110 26336
rect 16807 26268 17448 26296
rect 16807 26265 16819 26268
rect 16761 26259 16819 26265
rect 17678 26256 17684 26308
rect 17736 26256 17742 26308
rect 17773 26299 17831 26305
rect 17773 26265 17785 26299
rect 17819 26296 17831 26299
rect 18138 26296 18144 26308
rect 17819 26268 18144 26296
rect 17819 26265 17831 26268
rect 17773 26259 17831 26265
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 18248 26296 18276 26336
rect 18325 26333 18337 26367
rect 18371 26364 18383 26367
rect 18414 26364 18420 26376
rect 18371 26336 18420 26364
rect 18371 26333 18383 26336
rect 18325 26327 18383 26333
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18598 26324 18604 26376
rect 18656 26324 18662 26376
rect 18690 26324 18696 26376
rect 18748 26324 18754 26376
rect 18966 26324 18972 26376
rect 19024 26324 19030 26376
rect 19242 26324 19248 26376
rect 19300 26324 19306 26376
rect 18248 26268 18552 26296
rect 16390 26228 16396 26240
rect 16040 26200 16396 26228
rect 16390 26188 16396 26200
rect 16448 26228 16454 26240
rect 18417 26231 18475 26237
rect 18417 26228 18429 26231
rect 16448 26200 18429 26228
rect 16448 26188 16454 26200
rect 18417 26197 18429 26200
rect 18463 26197 18475 26231
rect 18524 26228 18552 26268
rect 18782 26256 18788 26308
rect 18840 26296 18846 26308
rect 19536 26296 19564 26404
rect 19610 26324 19616 26376
rect 19668 26324 19674 26376
rect 19812 26373 19840 26404
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20070 26364 20076 26376
rect 19843 26336 20076 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20070 26324 20076 26336
rect 20128 26364 20134 26376
rect 23201 26367 23259 26373
rect 20128 26336 20668 26364
rect 20128 26324 20134 26336
rect 18840 26268 19564 26296
rect 19628 26296 19656 26324
rect 19889 26299 19947 26305
rect 19889 26296 19901 26299
rect 19628 26268 19901 26296
rect 18840 26256 18846 26268
rect 19889 26265 19901 26268
rect 19935 26265 19947 26299
rect 19889 26259 19947 26265
rect 20254 26256 20260 26308
rect 20312 26296 20318 26308
rect 20349 26299 20407 26305
rect 20349 26296 20361 26299
rect 20312 26268 20361 26296
rect 20312 26256 20318 26268
rect 20349 26265 20361 26268
rect 20395 26265 20407 26299
rect 20349 26259 20407 26265
rect 19334 26228 19340 26240
rect 18524 26200 19340 26228
rect 18417 26191 18475 26197
rect 19334 26188 19340 26200
rect 19392 26188 19398 26240
rect 19794 26188 19800 26240
rect 19852 26228 19858 26240
rect 20549 26231 20607 26237
rect 20549 26228 20561 26231
rect 19852 26200 20561 26228
rect 19852 26188 19858 26200
rect 20549 26197 20561 26200
rect 20595 26197 20607 26231
rect 20640 26228 20668 26336
rect 23201 26333 23213 26367
rect 23247 26333 23259 26367
rect 23201 26327 23259 26333
rect 23293 26367 23351 26373
rect 23293 26333 23305 26367
rect 23339 26364 23351 26367
rect 23382 26364 23388 26376
rect 23339 26336 23388 26364
rect 23339 26333 23351 26336
rect 23293 26327 23351 26333
rect 23216 26296 23244 26327
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 23492 26364 23520 26463
rect 24762 26392 24768 26444
rect 24820 26432 24826 26444
rect 24949 26435 25007 26441
rect 24949 26432 24961 26435
rect 24820 26404 24961 26432
rect 24820 26392 24826 26404
rect 24949 26401 24961 26404
rect 24995 26401 25007 26435
rect 24949 26395 25007 26401
rect 25866 26392 25872 26444
rect 25924 26432 25930 26444
rect 26436 26432 26464 26472
rect 27433 26469 27445 26472
rect 27479 26469 27491 26503
rect 27433 26463 27491 26469
rect 27982 26460 27988 26512
rect 28040 26460 28046 26512
rect 25924 26404 26464 26432
rect 26697 26435 26755 26441
rect 25924 26392 25930 26404
rect 26697 26401 26709 26435
rect 26743 26432 26755 26435
rect 27249 26435 27307 26441
rect 27249 26432 27261 26435
rect 26743 26404 27261 26432
rect 26743 26401 26755 26404
rect 26697 26395 26755 26401
rect 27249 26401 27261 26404
rect 27295 26432 27307 26435
rect 27295 26404 27752 26432
rect 27295 26401 27307 26404
rect 27249 26395 27307 26401
rect 24029 26367 24087 26373
rect 24029 26364 24041 26367
rect 23492 26336 24041 26364
rect 24029 26333 24041 26336
rect 24075 26333 24087 26367
rect 24029 26327 24087 26333
rect 24213 26367 24271 26373
rect 24213 26333 24225 26367
rect 24259 26333 24271 26367
rect 24213 26327 24271 26333
rect 23216 26268 23428 26296
rect 21818 26228 21824 26240
rect 20640 26200 21824 26228
rect 20549 26191 20607 26197
rect 21818 26188 21824 26200
rect 21876 26188 21882 26240
rect 23400 26228 23428 26268
rect 23474 26256 23480 26308
rect 23532 26296 23538 26308
rect 23569 26299 23627 26305
rect 23569 26296 23581 26299
rect 23532 26268 23581 26296
rect 23532 26256 23538 26268
rect 23569 26265 23581 26268
rect 23615 26265 23627 26299
rect 23569 26259 23627 26265
rect 23658 26256 23664 26308
rect 23716 26296 23722 26308
rect 23769 26299 23827 26305
rect 23769 26296 23781 26299
rect 23716 26268 23781 26296
rect 23716 26256 23722 26268
rect 23769 26265 23781 26268
rect 23815 26265 23827 26299
rect 24228 26296 24256 26327
rect 26970 26324 26976 26376
rect 27028 26324 27034 26376
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26333 27123 26367
rect 27065 26327 27123 26333
rect 27157 26367 27215 26373
rect 27157 26333 27169 26367
rect 27203 26333 27215 26367
rect 27157 26327 27215 26333
rect 23769 26259 23827 26265
rect 23952 26268 24256 26296
rect 23676 26228 23704 26256
rect 23952 26240 23980 26268
rect 25222 26256 25228 26308
rect 25280 26256 25286 26308
rect 26234 26256 26240 26308
rect 26292 26256 26298 26308
rect 23400 26200 23704 26228
rect 23934 26188 23940 26240
rect 23992 26188 23998 26240
rect 26786 26188 26792 26240
rect 26844 26188 26850 26240
rect 27080 26228 27108 26327
rect 27172 26296 27200 26327
rect 27338 26324 27344 26376
rect 27396 26364 27402 26376
rect 27724 26373 27752 26404
rect 27617 26367 27675 26373
rect 27617 26364 27629 26367
rect 27396 26336 27629 26364
rect 27396 26324 27402 26336
rect 27617 26333 27629 26336
rect 27663 26333 27675 26367
rect 27617 26327 27675 26333
rect 27709 26367 27767 26373
rect 27709 26333 27721 26367
rect 27755 26333 27767 26367
rect 27709 26327 27767 26333
rect 28000 26296 28028 26460
rect 27172 26268 28028 26296
rect 29270 26256 29276 26308
rect 29328 26256 29334 26308
rect 27338 26228 27344 26240
rect 27080 26200 27344 26228
rect 27338 26188 27344 26200
rect 27396 26188 27402 26240
rect 27798 26188 27804 26240
rect 27856 26188 27862 26240
rect 1104 26138 29716 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 29716 26138
rect 1104 26064 29716 26086
rect 2590 25984 2596 26036
rect 2648 26024 2654 26036
rect 2648 25996 2774 26024
rect 2648 25984 2654 25996
rect 2746 25684 2774 25996
rect 5350 25984 5356 26036
rect 5408 26024 5414 26036
rect 5445 26027 5503 26033
rect 5445 26024 5457 26027
rect 5408 25996 5457 26024
rect 5408 25984 5414 25996
rect 5445 25993 5457 25996
rect 5491 25993 5503 26027
rect 5445 25987 5503 25993
rect 5994 25984 6000 26036
rect 6052 26024 6058 26036
rect 6181 26027 6239 26033
rect 6181 26024 6193 26027
rect 6052 25996 6193 26024
rect 6052 25984 6058 25996
rect 6181 25993 6193 25996
rect 6227 25993 6239 26027
rect 6181 25987 6239 25993
rect 6730 25984 6736 26036
rect 6788 26024 6794 26036
rect 10229 26027 10287 26033
rect 6788 25996 9352 26024
rect 6788 25984 6794 25996
rect 4706 25916 4712 25968
rect 4764 25916 4770 25968
rect 5813 25959 5871 25965
rect 5813 25925 5825 25959
rect 5859 25956 5871 25959
rect 6086 25956 6092 25968
rect 5859 25928 6092 25956
rect 5859 25925 5871 25928
rect 5813 25919 5871 25925
rect 6086 25916 6092 25928
rect 6144 25916 6150 25968
rect 8294 25956 8300 25968
rect 6196 25928 6684 25956
rect 3694 25848 3700 25900
rect 3752 25848 3758 25900
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25888 5687 25891
rect 5718 25888 5724 25900
rect 5675 25860 5724 25888
rect 5675 25857 5687 25860
rect 5629 25851 5687 25857
rect 5718 25848 5724 25860
rect 5776 25848 5782 25900
rect 5905 25891 5963 25897
rect 5905 25857 5917 25891
rect 5951 25857 5963 25891
rect 5905 25851 5963 25857
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25888 6055 25891
rect 6196 25888 6224 25928
rect 6656 25900 6684 25928
rect 6748 25928 8300 25956
rect 6043 25860 6224 25888
rect 6043 25857 6055 25860
rect 5997 25851 6055 25857
rect 3970 25780 3976 25832
rect 4028 25780 4034 25832
rect 5920 25820 5948 25851
rect 6270 25848 6276 25900
rect 6328 25888 6334 25900
rect 6457 25891 6515 25897
rect 6457 25888 6469 25891
rect 6328 25860 6469 25888
rect 6328 25848 6334 25860
rect 6457 25857 6469 25860
rect 6503 25857 6515 25891
rect 6457 25851 6515 25857
rect 6638 25848 6644 25900
rect 6696 25848 6702 25900
rect 6748 25829 6776 25928
rect 8294 25916 8300 25928
rect 8352 25956 8358 25968
rect 8352 25928 9076 25956
rect 8352 25916 8358 25928
rect 6914 25848 6920 25900
rect 6972 25888 6978 25900
rect 7009 25891 7067 25897
rect 7009 25888 7021 25891
rect 6972 25860 7021 25888
rect 6972 25848 6978 25860
rect 7009 25857 7021 25860
rect 7055 25857 7067 25891
rect 7009 25851 7067 25857
rect 7558 25848 7564 25900
rect 7616 25848 7622 25900
rect 7742 25897 7748 25900
rect 7709 25891 7748 25897
rect 7709 25857 7721 25891
rect 7709 25851 7748 25857
rect 7742 25848 7748 25851
rect 7800 25848 7806 25900
rect 7834 25848 7840 25900
rect 7892 25848 7898 25900
rect 7929 25891 7987 25897
rect 7929 25857 7941 25891
rect 7975 25857 7987 25891
rect 7929 25851 7987 25857
rect 8067 25891 8125 25897
rect 8067 25857 8079 25891
rect 8113 25888 8125 25891
rect 8389 25891 8447 25897
rect 8389 25888 8401 25891
rect 8113 25860 8401 25888
rect 8113 25857 8125 25860
rect 8067 25851 8125 25857
rect 8389 25857 8401 25860
rect 8435 25857 8447 25891
rect 8389 25851 8447 25857
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25857 8539 25891
rect 8481 25851 8539 25857
rect 8941 25891 8999 25897
rect 8941 25857 8953 25891
rect 8987 25857 8999 25891
rect 8941 25851 8999 25857
rect 6733 25823 6791 25829
rect 6733 25820 6745 25823
rect 5920 25792 6745 25820
rect 6733 25789 6745 25792
rect 6779 25789 6791 25823
rect 6733 25783 6791 25789
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 6546 25712 6552 25764
rect 6604 25752 6610 25764
rect 6840 25752 6868 25783
rect 7466 25780 7472 25832
rect 7524 25820 7530 25832
rect 7944 25820 7972 25851
rect 7524 25792 8432 25820
rect 7524 25780 7530 25792
rect 8404 25764 8432 25792
rect 6604 25724 6868 25752
rect 6604 25712 6610 25724
rect 7006 25712 7012 25764
rect 7064 25752 7070 25764
rect 8205 25755 8263 25761
rect 8205 25752 8217 25755
rect 7064 25724 8217 25752
rect 7064 25712 7070 25724
rect 8205 25721 8217 25724
rect 8251 25721 8263 25755
rect 8205 25715 8263 25721
rect 8386 25712 8392 25764
rect 8444 25712 8450 25764
rect 7098 25684 7104 25696
rect 2746 25656 7104 25684
rect 7098 25644 7104 25656
rect 7156 25644 7162 25696
rect 7193 25687 7251 25693
rect 7193 25653 7205 25687
rect 7239 25684 7251 25687
rect 7650 25684 7656 25696
rect 7239 25656 7656 25684
rect 7239 25653 7251 25656
rect 7193 25647 7251 25653
rect 7650 25644 7656 25656
rect 7708 25644 7714 25696
rect 7926 25644 7932 25696
rect 7984 25684 7990 25696
rect 8496 25684 8524 25851
rect 8956 25752 8984 25851
rect 9048 25829 9076 25928
rect 9214 25848 9220 25900
rect 9272 25848 9278 25900
rect 9324 25897 9352 25996
rect 10229 25993 10241 26027
rect 10275 26024 10287 26027
rect 10870 26024 10876 26036
rect 10275 25996 10876 26024
rect 10275 25993 10287 25996
rect 10229 25987 10287 25993
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 12434 26024 12440 26036
rect 11808 25996 12440 26024
rect 9600 25928 10456 25956
rect 9600 25897 9628 25928
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25857 9367 25891
rect 9309 25851 9367 25857
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25888 9551 25891
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 9539 25860 9597 25888
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 9585 25857 9597 25860
rect 9631 25857 9643 25891
rect 9585 25851 9643 25857
rect 9033 25823 9091 25829
rect 9033 25789 9045 25823
rect 9079 25789 9091 25823
rect 9324 25820 9352 25851
rect 9858 25848 9864 25900
rect 9916 25848 9922 25900
rect 10428 25897 10456 25928
rect 10413 25891 10471 25897
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25857 10839 25891
rect 10781 25851 10839 25857
rect 9766 25820 9772 25832
rect 9324 25792 9772 25820
rect 9033 25783 9091 25789
rect 9766 25780 9772 25792
rect 9824 25780 9830 25832
rect 9876 25820 9904 25848
rect 10597 25823 10655 25829
rect 10597 25820 10609 25823
rect 9876 25792 10609 25820
rect 10597 25789 10609 25792
rect 10643 25789 10655 25823
rect 10597 25783 10655 25789
rect 10686 25780 10692 25832
rect 10744 25780 10750 25832
rect 10796 25820 10824 25851
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 11808 25897 11836 25996
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 13541 26027 13599 26033
rect 13541 25993 13553 26027
rect 13587 26024 13599 26027
rect 13630 26024 13636 26036
rect 13587 25996 13636 26024
rect 13587 25993 13599 25996
rect 13541 25987 13599 25993
rect 13556 25956 13584 25987
rect 13630 25984 13636 25996
rect 13688 25984 13694 26036
rect 14369 26027 14427 26033
rect 14369 25993 14381 26027
rect 14415 26024 14427 26027
rect 14826 26024 14832 26036
rect 14415 25996 14832 26024
rect 14415 25993 14427 25996
rect 14369 25987 14427 25993
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 15194 25984 15200 26036
rect 15252 25984 15258 26036
rect 15746 26024 15752 26036
rect 15672 25996 15752 26024
rect 15010 25956 15016 25968
rect 12452 25928 13584 25956
rect 14752 25928 15016 25956
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 11020 25860 11529 25888
rect 11020 25848 11026 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11793 25891 11851 25897
rect 11793 25857 11805 25891
rect 11839 25857 11851 25891
rect 11793 25851 11851 25857
rect 11882 25848 11888 25900
rect 11940 25888 11946 25900
rect 11977 25891 12035 25897
rect 11977 25888 11989 25891
rect 11940 25860 11989 25888
rect 11940 25848 11946 25860
rect 11977 25857 11989 25860
rect 12023 25857 12035 25891
rect 11977 25851 12035 25857
rect 12250 25848 12256 25900
rect 12308 25848 12314 25900
rect 12452 25897 12480 25928
rect 12437 25891 12495 25897
rect 12437 25857 12449 25891
rect 12483 25857 12495 25891
rect 12437 25851 12495 25857
rect 12805 25891 12863 25897
rect 12805 25857 12817 25891
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 12820 25820 12848 25851
rect 12894 25848 12900 25900
rect 12952 25888 12958 25900
rect 13265 25891 13323 25897
rect 12952 25860 13124 25888
rect 12952 25848 12958 25860
rect 13096 25832 13124 25860
rect 13265 25857 13277 25891
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 10796 25792 12848 25820
rect 12989 25823 13047 25829
rect 9398 25752 9404 25764
rect 8956 25724 9404 25752
rect 9398 25712 9404 25724
rect 9456 25752 9462 25764
rect 9858 25752 9864 25764
rect 9456 25724 9864 25752
rect 9456 25712 9462 25724
rect 9858 25712 9864 25724
rect 9916 25712 9922 25764
rect 10137 25755 10195 25761
rect 10137 25721 10149 25755
rect 10183 25752 10195 25755
rect 10796 25752 10824 25792
rect 12989 25789 13001 25823
rect 13035 25789 13047 25823
rect 12989 25783 13047 25789
rect 12345 25755 12403 25761
rect 12345 25752 12357 25755
rect 10183 25724 10824 25752
rect 11992 25724 12357 25752
rect 10183 25721 10195 25724
rect 10137 25715 10195 25721
rect 7984 25656 8524 25684
rect 7984 25644 7990 25656
rect 9950 25644 9956 25696
rect 10008 25644 10014 25696
rect 11992 25693 12020 25724
rect 12345 25721 12357 25724
rect 12391 25721 12403 25755
rect 12345 25715 12403 25721
rect 12544 25724 12756 25752
rect 11977 25687 12035 25693
rect 11977 25653 11989 25687
rect 12023 25653 12035 25687
rect 11977 25647 12035 25653
rect 12161 25687 12219 25693
rect 12161 25653 12173 25687
rect 12207 25684 12219 25687
rect 12544 25684 12572 25724
rect 12207 25656 12572 25684
rect 12207 25653 12219 25656
rect 12161 25647 12219 25653
rect 12618 25644 12624 25696
rect 12676 25644 12682 25696
rect 12728 25684 12756 25724
rect 12802 25712 12808 25764
rect 12860 25752 12866 25764
rect 12897 25755 12955 25761
rect 12897 25752 12909 25755
rect 12860 25724 12909 25752
rect 12860 25712 12866 25724
rect 12897 25721 12909 25724
rect 12943 25721 12955 25755
rect 12897 25715 12955 25721
rect 13004 25684 13032 25783
rect 13078 25780 13084 25832
rect 13136 25780 13142 25832
rect 13280 25820 13308 25851
rect 13354 25848 13360 25900
rect 13412 25848 13418 25900
rect 13446 25848 13452 25900
rect 13504 25888 13510 25900
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 13504 25860 13645 25888
rect 13504 25848 13510 25860
rect 13633 25857 13645 25860
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 13906 25848 13912 25900
rect 13964 25888 13970 25900
rect 14093 25891 14151 25897
rect 14093 25888 14105 25891
rect 13964 25860 14105 25888
rect 13964 25848 13970 25860
rect 14093 25857 14105 25860
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 14550 25848 14556 25900
rect 14608 25848 14614 25900
rect 14752 25897 14780 25928
rect 15010 25916 15016 25928
rect 15068 25916 15074 25968
rect 15120 25928 15608 25956
rect 15120 25897 15148 25928
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25857 14979 25891
rect 14921 25851 14979 25857
rect 15105 25891 15163 25897
rect 15105 25857 15117 25891
rect 15151 25857 15163 25891
rect 15105 25851 15163 25857
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15473 25891 15531 25897
rect 15473 25857 15485 25891
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 13280 25792 13400 25820
rect 13372 25761 13400 25792
rect 14274 25780 14280 25832
rect 14332 25820 14338 25832
rect 14826 25820 14832 25832
rect 14332 25792 14832 25820
rect 14332 25780 14338 25792
rect 14826 25780 14832 25792
rect 14884 25780 14890 25832
rect 14936 25820 14964 25851
rect 15396 25820 15424 25851
rect 14936 25792 15424 25820
rect 13357 25755 13415 25761
rect 13357 25721 13369 25755
rect 13403 25721 13415 25755
rect 14936 25752 14964 25792
rect 13357 25715 13415 25721
rect 14476 25724 14964 25752
rect 14476 25696 14504 25724
rect 12728 25656 13032 25684
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13446 25684 13452 25696
rect 13228 25656 13452 25684
rect 13228 25644 13234 25656
rect 13446 25644 13452 25656
rect 13504 25644 13510 25696
rect 14185 25687 14243 25693
rect 14185 25653 14197 25687
rect 14231 25684 14243 25687
rect 14458 25684 14464 25696
rect 14231 25656 14464 25684
rect 14231 25653 14243 25656
rect 14185 25647 14243 25653
rect 14458 25644 14464 25656
rect 14516 25644 14522 25696
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 15488 25684 15516 25851
rect 15580 25820 15608 25928
rect 15672 25897 15700 25996
rect 15746 25984 15752 25996
rect 15804 25984 15810 26036
rect 15930 25984 15936 26036
rect 15988 25984 15994 26036
rect 16206 25984 16212 26036
rect 16264 26024 16270 26036
rect 17865 26027 17923 26033
rect 17865 26024 17877 26027
rect 16264 25996 17877 26024
rect 16264 25984 16270 25996
rect 17865 25993 17877 25996
rect 17911 25993 17923 26027
rect 17865 25987 17923 25993
rect 18598 25984 18604 26036
rect 18656 26024 18662 26036
rect 21637 26027 21695 26033
rect 21637 26024 21649 26027
rect 18656 25996 21649 26024
rect 18656 25984 18662 25996
rect 16669 25959 16727 25965
rect 16669 25956 16681 25959
rect 15764 25928 16681 25956
rect 15764 25897 15792 25928
rect 16669 25925 16681 25928
rect 16715 25925 16727 25959
rect 16669 25919 16727 25925
rect 17034 25916 17040 25968
rect 17092 25956 17098 25968
rect 17678 25956 17684 25968
rect 17092 25928 17684 25956
rect 17092 25916 17098 25928
rect 17678 25916 17684 25928
rect 17736 25956 17742 25968
rect 18966 25956 18972 25968
rect 17736 25928 17908 25956
rect 17736 25916 17742 25928
rect 17880 25900 17908 25928
rect 18432 25928 18972 25956
rect 18432 25900 18460 25928
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25857 15715 25891
rect 15657 25851 15715 25857
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 15838 25848 15844 25900
rect 15896 25888 15902 25900
rect 16117 25891 16175 25897
rect 16117 25888 16129 25891
rect 15896 25860 16129 25888
rect 15896 25848 15902 25860
rect 16117 25857 16129 25860
rect 16163 25857 16175 25891
rect 16117 25851 16175 25857
rect 16485 25891 16543 25897
rect 16485 25857 16497 25891
rect 16531 25857 16543 25891
rect 16485 25851 16543 25857
rect 16206 25820 16212 25832
rect 15580 25792 16212 25820
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 16500 25820 16528 25851
rect 16850 25848 16856 25900
rect 16908 25848 16914 25900
rect 17126 25848 17132 25900
rect 17184 25848 17190 25900
rect 17862 25848 17868 25900
rect 17920 25848 17926 25900
rect 18046 25848 18052 25900
rect 18104 25848 18110 25900
rect 18138 25848 18144 25900
rect 18196 25848 18202 25900
rect 18414 25848 18420 25900
rect 18472 25848 18478 25900
rect 19260 25897 19288 25996
rect 21637 25993 21649 25996
rect 21683 25993 21695 26027
rect 21637 25987 21695 25993
rect 21818 25984 21824 26036
rect 21876 25984 21882 26036
rect 24486 25984 24492 26036
rect 24544 26024 24550 26036
rect 24765 26027 24823 26033
rect 24765 26024 24777 26027
rect 24544 25996 24777 26024
rect 24544 25984 24550 25996
rect 24765 25993 24777 25996
rect 24811 25993 24823 26027
rect 24765 25987 24823 25993
rect 25222 25984 25228 26036
rect 25280 26024 25286 26036
rect 25501 26027 25559 26033
rect 25501 26024 25513 26027
rect 25280 25996 25513 26024
rect 25280 25984 25286 25996
rect 25501 25993 25513 25996
rect 25547 25993 25559 26027
rect 25501 25987 25559 25993
rect 26145 26027 26203 26033
rect 26145 25993 26157 26027
rect 26191 26024 26203 26027
rect 26234 26024 26240 26036
rect 26191 25996 26240 26024
rect 26191 25993 26203 25996
rect 26145 25987 26203 25993
rect 26234 25984 26240 25996
rect 26292 25984 26298 26036
rect 27798 26024 27804 26036
rect 27356 25996 27804 26024
rect 27356 25968 27384 25996
rect 27798 25984 27804 25996
rect 27856 26024 27862 26036
rect 29365 26027 29423 26033
rect 29365 26024 29377 26027
rect 27856 25996 29377 26024
rect 27856 25984 27862 25996
rect 29365 25993 29377 25996
rect 29411 25993 29423 26027
rect 29365 25987 29423 25993
rect 19426 25956 19432 25968
rect 19352 25928 19432 25956
rect 19352 25897 19380 25928
rect 19426 25916 19432 25928
rect 19484 25956 19490 25968
rect 20254 25956 20260 25968
rect 19484 25928 20260 25956
rect 19484 25916 19490 25928
rect 20254 25916 20260 25928
rect 20312 25916 20318 25968
rect 21450 25956 21456 25968
rect 21390 25928 21456 25956
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 22278 25916 22284 25968
rect 22336 25916 22342 25968
rect 23290 25916 23296 25968
rect 23348 25916 23354 25968
rect 25866 25916 25872 25968
rect 25924 25956 25930 25968
rect 25961 25959 26019 25965
rect 25961 25956 25973 25959
rect 25924 25928 25973 25956
rect 25924 25916 25930 25928
rect 25961 25925 25973 25928
rect 26007 25925 26019 25959
rect 25961 25919 26019 25925
rect 27338 25916 27344 25968
rect 27396 25916 27402 25968
rect 18509 25891 18567 25897
rect 18509 25857 18521 25891
rect 18555 25888 18567 25891
rect 19245 25891 19303 25897
rect 18555 25860 18920 25888
rect 18555 25857 18567 25860
rect 18509 25851 18567 25857
rect 17586 25820 17592 25832
rect 16500 25792 17592 25820
rect 17586 25780 17592 25792
rect 17644 25780 17650 25832
rect 18156 25820 18184 25848
rect 18601 25823 18659 25829
rect 18601 25820 18613 25823
rect 18156 25792 18613 25820
rect 18601 25789 18613 25792
rect 18647 25789 18659 25823
rect 18601 25783 18659 25789
rect 18325 25755 18383 25761
rect 18325 25721 18337 25755
rect 18371 25752 18383 25755
rect 18782 25752 18788 25764
rect 18371 25724 18788 25752
rect 18371 25721 18383 25724
rect 18325 25715 18383 25721
rect 18782 25712 18788 25724
rect 18840 25712 18846 25764
rect 14884 25656 15516 25684
rect 14884 25644 14890 25656
rect 16390 25644 16396 25696
rect 16448 25644 16454 25696
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 18892 25684 18920 25860
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 19337 25891 19395 25897
rect 19337 25857 19349 25891
rect 19383 25857 19395 25891
rect 19705 25891 19763 25897
rect 19705 25888 19717 25891
rect 19337 25851 19395 25857
rect 19444 25860 19717 25888
rect 19444 25764 19472 25860
rect 19705 25857 19717 25860
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 19794 25848 19800 25900
rect 19852 25848 19858 25900
rect 19886 25848 19892 25900
rect 19944 25848 19950 25900
rect 23569 25891 23627 25897
rect 23569 25857 23581 25891
rect 23615 25888 23627 25891
rect 24762 25888 24768 25900
rect 23615 25860 24768 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 24762 25848 24768 25860
rect 24820 25848 24826 25900
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25888 24915 25891
rect 26234 25888 26240 25900
rect 24903 25860 26240 25888
rect 24903 25857 24915 25860
rect 24857 25851 24915 25857
rect 19521 25823 19579 25829
rect 19521 25789 19533 25823
rect 19567 25820 19579 25823
rect 20165 25823 20223 25829
rect 20165 25820 20177 25823
rect 19567 25792 20177 25820
rect 19567 25789 19579 25792
rect 19521 25783 19579 25789
rect 20165 25789 20177 25792
rect 20211 25789 20223 25823
rect 20165 25783 20223 25789
rect 22002 25780 22008 25832
rect 22060 25820 22066 25832
rect 24872 25820 24900 25851
rect 26234 25848 26240 25860
rect 26292 25848 26298 25900
rect 27154 25848 27160 25900
rect 27212 25848 27218 25900
rect 28994 25848 29000 25900
rect 29052 25848 29058 25900
rect 22060 25792 24900 25820
rect 22060 25780 22066 25792
rect 27614 25780 27620 25832
rect 27672 25780 27678 25832
rect 27893 25823 27951 25829
rect 27893 25789 27905 25823
rect 27939 25820 27951 25823
rect 27982 25820 27988 25832
rect 27939 25792 27988 25820
rect 27939 25789 27951 25792
rect 27893 25783 27951 25789
rect 27982 25780 27988 25792
rect 28040 25780 28046 25832
rect 19153 25755 19211 25761
rect 19153 25721 19165 25755
rect 19199 25752 19211 25755
rect 19426 25752 19432 25764
rect 19199 25724 19432 25752
rect 19199 25721 19211 25724
rect 19153 25715 19211 25721
rect 19426 25712 19432 25724
rect 19484 25712 19490 25764
rect 25685 25755 25743 25761
rect 25685 25721 25697 25755
rect 25731 25752 25743 25755
rect 26786 25752 26792 25764
rect 25731 25724 26792 25752
rect 25731 25721 25743 25724
rect 25685 25715 25743 25721
rect 26786 25712 26792 25724
rect 26844 25712 26850 25764
rect 17460 25656 18920 25684
rect 27525 25687 27583 25693
rect 17460 25644 17466 25656
rect 27525 25653 27537 25687
rect 27571 25684 27583 25687
rect 27706 25684 27712 25696
rect 27571 25656 27712 25684
rect 27571 25653 27583 25656
rect 27525 25647 27583 25653
rect 27706 25644 27712 25656
rect 27764 25644 27770 25696
rect 1104 25594 29716 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 29716 25594
rect 1104 25520 29716 25542
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 4157 25483 4215 25489
rect 4157 25480 4169 25483
rect 4028 25452 4169 25480
rect 4028 25440 4034 25452
rect 4157 25449 4169 25452
rect 4203 25449 4215 25483
rect 4157 25443 4215 25449
rect 4341 25483 4399 25489
rect 4341 25449 4353 25483
rect 4387 25480 4399 25483
rect 4614 25480 4620 25492
rect 4387 25452 4620 25480
rect 4387 25449 4399 25452
rect 4341 25443 4399 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 9214 25440 9220 25492
rect 9272 25480 9278 25492
rect 9674 25480 9680 25492
rect 9272 25452 9680 25480
rect 9272 25440 9278 25452
rect 9674 25440 9680 25452
rect 9732 25440 9738 25492
rect 9950 25440 9956 25492
rect 10008 25440 10014 25492
rect 11882 25440 11888 25492
rect 11940 25440 11946 25492
rect 12897 25483 12955 25489
rect 12897 25449 12909 25483
rect 12943 25480 12955 25483
rect 12986 25480 12992 25492
rect 12943 25452 12992 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 12986 25440 12992 25452
rect 13044 25480 13050 25492
rect 13354 25480 13360 25492
rect 13044 25452 13360 25480
rect 13044 25440 13050 25452
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 14458 25440 14464 25492
rect 14516 25440 14522 25492
rect 16301 25483 16359 25489
rect 16301 25449 16313 25483
rect 16347 25480 16359 25483
rect 16942 25480 16948 25492
rect 16347 25452 16948 25480
rect 16347 25449 16359 25452
rect 16301 25443 16359 25449
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 17586 25440 17592 25492
rect 17644 25440 17650 25492
rect 18414 25440 18420 25492
rect 18472 25480 18478 25492
rect 18509 25483 18567 25489
rect 18509 25480 18521 25483
rect 18472 25452 18521 25480
rect 18472 25440 18478 25452
rect 18509 25449 18521 25452
rect 18555 25449 18567 25483
rect 18509 25443 18567 25449
rect 21450 25440 21456 25492
rect 21508 25440 21514 25492
rect 22278 25440 22284 25492
rect 22336 25440 22342 25492
rect 27341 25483 27399 25489
rect 27341 25449 27353 25483
rect 27387 25480 27399 25483
rect 27430 25480 27436 25492
rect 27387 25452 27436 25480
rect 27387 25449 27399 25452
rect 27341 25443 27399 25449
rect 27430 25440 27436 25452
rect 27488 25440 27494 25492
rect 27982 25440 27988 25492
rect 28040 25440 28046 25492
rect 28813 25483 28871 25489
rect 28813 25449 28825 25483
rect 28859 25480 28871 25483
rect 28994 25480 29000 25492
rect 28859 25452 29000 25480
rect 28859 25449 28871 25452
rect 28813 25443 28871 25449
rect 28994 25440 29000 25452
rect 29052 25440 29058 25492
rect 6270 25372 6276 25424
rect 6328 25412 6334 25424
rect 7837 25415 7895 25421
rect 6328 25384 7696 25412
rect 6328 25372 6334 25384
rect 7101 25347 7159 25353
rect 7101 25313 7113 25347
rect 7147 25344 7159 25347
rect 7668 25344 7696 25384
rect 7837 25381 7849 25415
rect 7883 25412 7895 25415
rect 7926 25412 7932 25424
rect 7883 25384 7932 25412
rect 7883 25381 7895 25384
rect 7837 25375 7895 25381
rect 7926 25372 7932 25384
rect 7984 25372 7990 25424
rect 10686 25372 10692 25424
rect 10744 25412 10750 25424
rect 11333 25415 11391 25421
rect 11333 25412 11345 25415
rect 10744 25384 11345 25412
rect 10744 25372 10750 25384
rect 11333 25381 11345 25384
rect 11379 25412 11391 25415
rect 12250 25412 12256 25424
rect 11379 25384 12256 25412
rect 11379 25381 11391 25384
rect 11333 25375 11391 25381
rect 12250 25372 12256 25384
rect 12308 25372 12314 25424
rect 13078 25372 13084 25424
rect 13136 25412 13142 25424
rect 13541 25415 13599 25421
rect 13541 25412 13553 25415
rect 13136 25384 13553 25412
rect 13136 25372 13142 25384
rect 13541 25381 13553 25384
rect 13587 25381 13599 25415
rect 13541 25375 13599 25381
rect 17034 25372 17040 25424
rect 17092 25412 17098 25424
rect 17092 25384 17172 25412
rect 17092 25372 17098 25384
rect 7147 25316 7604 25344
rect 7668 25316 8248 25344
rect 7147 25313 7159 25316
rect 7101 25307 7159 25313
rect 7576 25288 7604 25316
rect 4706 25236 4712 25288
rect 4764 25276 4770 25288
rect 5902 25276 5908 25288
rect 4764 25248 5908 25276
rect 4764 25236 4770 25248
rect 5902 25236 5908 25248
rect 5960 25236 5966 25288
rect 5994 25236 6000 25288
rect 6052 25276 6058 25288
rect 6362 25285 6368 25288
rect 6181 25279 6239 25285
rect 6181 25276 6193 25279
rect 6052 25248 6193 25276
rect 6052 25236 6058 25248
rect 6181 25245 6193 25248
rect 6227 25245 6239 25279
rect 6181 25239 6239 25245
rect 6329 25279 6368 25285
rect 6329 25245 6341 25279
rect 6329 25239 6368 25245
rect 6362 25236 6368 25239
rect 6420 25236 6426 25288
rect 6730 25285 6736 25288
rect 6687 25279 6736 25285
rect 6687 25276 6699 25279
rect 6643 25248 6699 25276
rect 6687 25245 6699 25248
rect 6733 25245 6736 25279
rect 6687 25239 6736 25245
rect 6730 25236 6736 25239
rect 6788 25276 6794 25288
rect 7009 25279 7067 25285
rect 7009 25276 7021 25279
rect 6788 25248 7021 25276
rect 6788 25236 6794 25248
rect 7009 25245 7021 25248
rect 7055 25245 7067 25279
rect 7009 25239 7067 25245
rect 7190 25236 7196 25288
rect 7248 25236 7254 25288
rect 7558 25236 7564 25288
rect 7616 25236 7622 25288
rect 7650 25236 7656 25288
rect 7708 25236 7714 25288
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25276 7987 25279
rect 7975 25248 8156 25276
rect 7975 25245 7987 25248
rect 7929 25239 7987 25245
rect 6454 25168 6460 25220
rect 6512 25168 6518 25220
rect 6549 25211 6607 25217
rect 6549 25177 6561 25211
rect 6595 25208 6607 25211
rect 7208 25208 7236 25236
rect 8018 25208 8024 25220
rect 6595 25180 8024 25208
rect 6595 25177 6607 25180
rect 6549 25171 6607 25177
rect 8018 25168 8024 25180
rect 8076 25168 8082 25220
rect 8128 25152 8156 25248
rect 8220 25208 8248 25316
rect 8386 25304 8392 25356
rect 8444 25344 8450 25356
rect 10873 25347 10931 25353
rect 8444 25316 8708 25344
rect 8444 25304 8450 25316
rect 8680 25288 8708 25316
rect 9416 25316 10824 25344
rect 8662 25236 8668 25288
rect 8720 25236 8726 25288
rect 9416 25285 9444 25316
rect 9401 25279 9459 25285
rect 9401 25245 9413 25279
rect 9447 25245 9459 25279
rect 9401 25239 9459 25245
rect 9674 25236 9680 25288
rect 9732 25236 9738 25288
rect 9766 25236 9772 25288
rect 9824 25276 9830 25288
rect 10594 25276 10600 25288
rect 9824 25248 10600 25276
rect 9824 25236 9830 25248
rect 10594 25236 10600 25248
rect 10652 25236 10658 25288
rect 10686 25236 10692 25288
rect 10744 25276 10750 25288
rect 10796 25285 10824 25316
rect 10873 25313 10885 25347
rect 10919 25313 10931 25347
rect 10873 25307 10931 25313
rect 10781 25279 10839 25285
rect 10781 25276 10793 25279
rect 10744 25248 10793 25276
rect 10744 25236 10750 25248
rect 10781 25245 10793 25248
rect 10827 25245 10839 25279
rect 10781 25239 10839 25245
rect 9585 25211 9643 25217
rect 9585 25208 9597 25211
rect 8220 25180 9597 25208
rect 9585 25177 9597 25180
rect 9631 25208 9643 25211
rect 10410 25208 10416 25220
rect 9631 25180 10416 25208
rect 9631 25177 9643 25180
rect 9585 25171 9643 25177
rect 10410 25168 10416 25180
rect 10468 25208 10474 25220
rect 10888 25208 10916 25307
rect 11238 25304 11244 25356
rect 11296 25344 11302 25356
rect 13262 25344 13268 25356
rect 11296 25316 11744 25344
rect 11296 25304 11302 25316
rect 11057 25279 11115 25285
rect 11057 25245 11069 25279
rect 11103 25245 11115 25279
rect 11057 25239 11115 25245
rect 10468 25180 10916 25208
rect 11072 25208 11100 25239
rect 11146 25236 11152 25288
rect 11204 25276 11210 25288
rect 11716 25285 11744 25316
rect 13096 25316 13268 25344
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11204 25248 11437 25276
rect 11204 25236 11210 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11701 25279 11759 25285
rect 11701 25245 11713 25279
rect 11747 25245 11759 25279
rect 11701 25239 11759 25245
rect 12894 25236 12900 25288
rect 12952 25276 12958 25288
rect 13096 25285 13124 25316
rect 13262 25304 13268 25316
rect 13320 25344 13326 25356
rect 17144 25353 17172 25384
rect 14645 25347 14703 25353
rect 13320 25316 13584 25344
rect 13320 25304 13326 25316
rect 13081 25279 13139 25285
rect 13081 25276 13093 25279
rect 12952 25248 13093 25276
rect 12952 25236 12958 25248
rect 13081 25245 13093 25248
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 13446 25236 13452 25288
rect 13504 25236 13510 25288
rect 13556 25285 13584 25316
rect 14645 25313 14657 25347
rect 14691 25344 14703 25347
rect 15933 25347 15991 25353
rect 15933 25344 15945 25347
rect 14691 25316 15945 25344
rect 14691 25313 14703 25316
rect 14645 25307 14703 25313
rect 15933 25313 15945 25316
rect 15979 25313 15991 25347
rect 15933 25307 15991 25313
rect 17129 25347 17187 25353
rect 17129 25313 17141 25347
rect 17175 25313 17187 25347
rect 17129 25307 17187 25313
rect 17221 25347 17279 25353
rect 17221 25313 17233 25347
rect 17267 25344 17279 25347
rect 17862 25344 17868 25356
rect 17267 25316 17868 25344
rect 17267 25313 17279 25316
rect 17221 25307 17279 25313
rect 17862 25304 17868 25316
rect 17920 25344 17926 25356
rect 19702 25344 19708 25356
rect 17920 25316 19708 25344
rect 17920 25304 17926 25316
rect 19702 25304 19708 25316
rect 19760 25344 19766 25356
rect 20530 25344 20536 25356
rect 19760 25316 20536 25344
rect 19760 25304 19766 25316
rect 20530 25304 20536 25316
rect 20588 25304 20594 25356
rect 27448 25344 27476 25440
rect 27617 25347 27675 25353
rect 27617 25344 27629 25347
rect 27448 25316 27629 25344
rect 27617 25313 27629 25316
rect 27663 25313 27675 25347
rect 27617 25307 27675 25313
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25245 13599 25279
rect 13541 25239 13599 25245
rect 13725 25279 13783 25285
rect 13725 25245 13737 25279
rect 13771 25245 13783 25279
rect 13725 25239 13783 25245
rect 11072 25180 11560 25208
rect 10468 25168 10474 25180
rect 3878 25100 3884 25152
rect 3936 25140 3942 25152
rect 4341 25143 4399 25149
rect 4341 25140 4353 25143
rect 3936 25112 4353 25140
rect 3936 25100 3942 25112
rect 4341 25109 4353 25112
rect 4387 25140 4399 25143
rect 6178 25140 6184 25152
rect 4387 25112 6184 25140
rect 4387 25109 4399 25112
rect 4341 25103 4399 25109
rect 6178 25100 6184 25112
rect 6236 25100 6242 25152
rect 6822 25100 6828 25152
rect 6880 25100 6886 25152
rect 7374 25100 7380 25152
rect 7432 25100 7438 25152
rect 8110 25100 8116 25152
rect 8168 25140 8174 25152
rect 8573 25143 8631 25149
rect 8573 25140 8585 25143
rect 8168 25112 8585 25140
rect 8168 25100 8174 25112
rect 8573 25109 8585 25112
rect 8619 25140 8631 25143
rect 9766 25140 9772 25152
rect 8619 25112 9772 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 9766 25100 9772 25112
rect 9824 25100 9830 25152
rect 11532 25149 11560 25180
rect 13170 25168 13176 25220
rect 13228 25168 13234 25220
rect 13262 25168 13268 25220
rect 13320 25208 13326 25220
rect 13630 25208 13636 25220
rect 13320 25180 13636 25208
rect 13320 25168 13326 25180
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 11517 25143 11575 25149
rect 11517 25109 11529 25143
rect 11563 25140 11575 25143
rect 12342 25140 12348 25152
rect 11563 25112 12348 25140
rect 11563 25109 11575 25112
rect 11517 25103 11575 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 13188 25140 13216 25168
rect 13740 25140 13768 25239
rect 14274 25236 14280 25288
rect 14332 25276 14338 25288
rect 14553 25279 14611 25285
rect 14553 25276 14565 25279
rect 14332 25248 14565 25276
rect 14332 25236 14338 25248
rect 14553 25245 14565 25248
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 15838 25236 15844 25288
rect 15896 25236 15902 25288
rect 16117 25279 16175 25285
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16666 25276 16672 25288
rect 16163 25248 16672 25276
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16666 25236 16672 25248
rect 16724 25276 16730 25288
rect 16853 25279 16911 25285
rect 16853 25276 16865 25279
rect 16724 25248 16865 25276
rect 16724 25236 16730 25248
rect 16853 25245 16865 25248
rect 16899 25245 16911 25279
rect 16853 25239 16911 25245
rect 17034 25236 17040 25288
rect 17092 25236 17098 25288
rect 17402 25236 17408 25288
rect 17460 25236 17466 25288
rect 18506 25236 18512 25288
rect 18564 25276 18570 25288
rect 18601 25279 18659 25285
rect 18601 25276 18613 25279
rect 18564 25248 18613 25276
rect 18564 25236 18570 25248
rect 18601 25245 18613 25248
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20070 25276 20076 25288
rect 19935 25248 20076 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25276 21603 25279
rect 22002 25276 22008 25288
rect 21591 25248 22008 25276
rect 21591 25245 21603 25248
rect 21545 25239 21603 25245
rect 22002 25236 22008 25248
rect 22060 25276 22066 25288
rect 22189 25279 22247 25285
rect 22189 25276 22201 25279
rect 22060 25248 22201 25276
rect 22060 25236 22066 25248
rect 22189 25245 22201 25248
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25276 23443 25279
rect 23566 25276 23572 25288
rect 23431 25248 23572 25276
rect 23431 25245 23443 25248
rect 23385 25239 23443 25245
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 23661 25279 23719 25285
rect 23661 25245 23673 25279
rect 23707 25276 23719 25279
rect 23750 25276 23756 25288
rect 23707 25248 23756 25276
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 26786 25236 26792 25288
rect 26844 25276 26850 25288
rect 27154 25276 27160 25288
rect 26844 25248 27160 25276
rect 26844 25236 26850 25248
rect 27154 25236 27160 25248
rect 27212 25276 27218 25288
rect 27249 25279 27307 25285
rect 27249 25276 27261 25279
rect 27212 25248 27261 25276
rect 27212 25236 27218 25248
rect 27249 25245 27261 25248
rect 27295 25245 27307 25279
rect 27249 25239 27307 25245
rect 27338 25236 27344 25288
rect 27396 25276 27402 25288
rect 27433 25279 27491 25285
rect 27433 25276 27445 25279
rect 27396 25248 27445 25276
rect 27396 25236 27402 25248
rect 27433 25245 27445 25248
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 27706 25236 27712 25288
rect 27764 25276 27770 25288
rect 27801 25279 27859 25285
rect 27801 25276 27813 25279
rect 27764 25248 27813 25276
rect 27764 25236 27770 25248
rect 27801 25245 27813 25248
rect 27847 25245 27859 25279
rect 27801 25239 27859 25245
rect 28905 25279 28963 25285
rect 28905 25245 28917 25279
rect 28951 25276 28963 25279
rect 29086 25276 29092 25288
rect 28951 25248 29092 25276
rect 28951 25245 28963 25248
rect 28905 25239 28963 25245
rect 14182 25168 14188 25220
rect 14240 25168 14246 25220
rect 26234 25168 26240 25220
rect 26292 25208 26298 25220
rect 28920 25208 28948 25239
rect 29086 25236 29092 25248
rect 29144 25236 29150 25288
rect 26292 25180 28948 25208
rect 26292 25168 26298 25180
rect 13188 25112 13768 25140
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14642 25140 14648 25152
rect 14323 25112 14648 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14642 25100 14648 25112
rect 14700 25100 14706 25152
rect 15930 25100 15936 25152
rect 15988 25140 15994 25152
rect 19518 25140 19524 25152
rect 15988 25112 19524 25140
rect 15988 25100 15994 25112
rect 19518 25100 19524 25112
rect 19576 25100 19582 25152
rect 19794 25100 19800 25152
rect 19852 25100 19858 25152
rect 23106 25100 23112 25152
rect 23164 25140 23170 25152
rect 23201 25143 23259 25149
rect 23201 25140 23213 25143
rect 23164 25112 23213 25140
rect 23164 25100 23170 25112
rect 23201 25109 23213 25112
rect 23247 25109 23259 25143
rect 23201 25103 23259 25109
rect 23569 25143 23627 25149
rect 23569 25109 23581 25143
rect 23615 25140 23627 25143
rect 24026 25140 24032 25152
rect 23615 25112 24032 25140
rect 23615 25109 23627 25112
rect 23569 25103 23627 25109
rect 24026 25100 24032 25112
rect 24084 25100 24090 25152
rect 1104 25050 29716 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 29716 25050
rect 1104 24976 29716 24998
rect 5166 24896 5172 24948
rect 5224 24936 5230 24948
rect 5350 24936 5356 24948
rect 5224 24908 5356 24936
rect 5224 24896 5230 24908
rect 5350 24896 5356 24908
rect 5408 24896 5414 24948
rect 5626 24896 5632 24948
rect 5684 24896 5690 24948
rect 5902 24896 5908 24948
rect 5960 24936 5966 24948
rect 6641 24939 6699 24945
rect 6641 24936 6653 24939
rect 5960 24908 6653 24936
rect 5960 24896 5966 24908
rect 6641 24905 6653 24908
rect 6687 24905 6699 24939
rect 6641 24899 6699 24905
rect 6822 24896 6828 24948
rect 6880 24896 6886 24948
rect 7098 24896 7104 24948
rect 7156 24936 7162 24948
rect 14274 24936 14280 24948
rect 7156 24908 14280 24936
rect 7156 24896 7162 24908
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 15749 24939 15807 24945
rect 15749 24905 15761 24939
rect 15795 24936 15807 24939
rect 15838 24936 15844 24948
rect 15795 24908 15844 24936
rect 15795 24905 15807 24908
rect 15749 24899 15807 24905
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 16666 24896 16672 24948
rect 16724 24896 16730 24948
rect 16850 24896 16856 24948
rect 16908 24936 16914 24948
rect 17405 24939 17463 24945
rect 17405 24936 17417 24939
rect 16908 24908 17417 24936
rect 16908 24896 16914 24908
rect 17405 24905 17417 24908
rect 17451 24905 17463 24939
rect 21266 24936 21272 24948
rect 17405 24899 17463 24905
rect 18064 24908 21272 24936
rect 6840 24868 6868 24896
rect 6840 24840 6960 24868
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 5350 24760 5356 24812
rect 5408 24800 5414 24812
rect 5570 24803 5628 24809
rect 5570 24800 5582 24803
rect 5408 24772 5582 24800
rect 5408 24760 5414 24772
rect 5570 24769 5582 24772
rect 5616 24769 5628 24803
rect 5570 24763 5628 24769
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 6089 24803 6147 24809
rect 6089 24800 6101 24803
rect 5776 24772 6101 24800
rect 5776 24760 5782 24772
rect 6089 24769 6101 24772
rect 6135 24800 6147 24803
rect 6638 24800 6644 24812
rect 6135 24772 6644 24800
rect 6135 24769 6147 24772
rect 6089 24763 6147 24769
rect 6638 24760 6644 24772
rect 6696 24760 6702 24812
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24769 6883 24803
rect 6932 24800 6960 24840
rect 7374 24828 7380 24880
rect 7432 24868 7438 24880
rect 7745 24871 7803 24877
rect 7745 24868 7757 24871
rect 7432 24840 7757 24868
rect 7432 24828 7438 24840
rect 7745 24837 7757 24840
rect 7791 24837 7803 24871
rect 7745 24831 7803 24837
rect 7834 24828 7840 24880
rect 7892 24868 7898 24880
rect 7892 24840 8064 24868
rect 7892 24828 7898 24840
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 6932 24772 7113 24800
rect 6825 24763 6883 24769
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7929 24803 7987 24809
rect 7929 24800 7941 24803
rect 7101 24763 7159 24769
rect 7484 24772 7941 24800
rect 5258 24624 5264 24676
rect 5316 24664 5322 24676
rect 5445 24667 5503 24673
rect 5445 24664 5457 24667
rect 5316 24636 5457 24664
rect 5316 24624 5322 24636
rect 5445 24633 5457 24636
rect 5491 24633 5503 24667
rect 5445 24627 5503 24633
rect 5626 24624 5632 24676
rect 5684 24664 5690 24676
rect 6840 24664 6868 24763
rect 7006 24692 7012 24744
rect 7064 24692 7070 24744
rect 7484 24664 7512 24772
rect 7929 24769 7941 24772
rect 7975 24769 7987 24803
rect 8036 24800 8064 24840
rect 8662 24828 8668 24880
rect 8720 24868 8726 24880
rect 9582 24868 9588 24880
rect 8720 24840 9588 24868
rect 8720 24828 8726 24840
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 15930 24868 15936 24880
rect 9692 24840 15936 24868
rect 9692 24800 9720 24840
rect 15930 24828 15936 24840
rect 15988 24828 15994 24880
rect 17954 24868 17960 24880
rect 16868 24840 17960 24868
rect 8036 24772 9720 24800
rect 7929 24763 7987 24769
rect 10042 24760 10048 24812
rect 10100 24760 10106 24812
rect 10502 24760 10508 24812
rect 10560 24800 10566 24812
rect 10560 24772 12388 24800
rect 10560 24760 10566 24772
rect 8662 24692 8668 24744
rect 8720 24732 8726 24744
rect 12250 24732 12256 24744
rect 8720 24704 12256 24732
rect 8720 24692 8726 24704
rect 12250 24692 12256 24704
rect 12308 24692 12314 24744
rect 12360 24732 12388 24772
rect 14642 24760 14648 24812
rect 14700 24760 14706 24812
rect 14734 24760 14740 24812
rect 14792 24800 14798 24812
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 14792 24772 15209 24800
rect 14792 24760 14798 24772
rect 15197 24769 15209 24772
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 15378 24760 15384 24812
rect 15436 24760 15442 24812
rect 15470 24760 15476 24812
rect 15528 24760 15534 24812
rect 15562 24760 15568 24812
rect 15620 24800 15626 24812
rect 16868 24809 16896 24840
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 15620 24772 16865 24800
rect 15620 24760 15626 24772
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 16942 24760 16948 24812
rect 17000 24760 17006 24812
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 17184 24772 17233 24800
rect 17184 24760 17190 24772
rect 17221 24769 17233 24772
rect 17267 24769 17279 24803
rect 17221 24763 17279 24769
rect 17310 24760 17316 24812
rect 17368 24760 17374 24812
rect 17494 24760 17500 24812
rect 17552 24760 17558 24812
rect 17589 24803 17647 24809
rect 17589 24769 17601 24803
rect 17635 24800 17647 24803
rect 17770 24800 17776 24812
rect 17635 24772 17776 24800
rect 17635 24769 17647 24772
rect 17589 24763 17647 24769
rect 17770 24760 17776 24772
rect 17828 24800 17834 24812
rect 18064 24800 18092 24908
rect 21266 24896 21272 24908
rect 21324 24896 21330 24948
rect 24121 24939 24179 24945
rect 24121 24905 24133 24939
rect 24167 24905 24179 24939
rect 24121 24899 24179 24905
rect 20070 24868 20076 24880
rect 19812 24840 20076 24868
rect 17828 24772 18092 24800
rect 17828 24760 17834 24772
rect 18414 24760 18420 24812
rect 18472 24800 18478 24812
rect 18693 24803 18751 24809
rect 18693 24800 18705 24803
rect 18472 24772 18705 24800
rect 18472 24760 18478 24772
rect 18693 24769 18705 24772
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 18874 24760 18880 24812
rect 18932 24760 18938 24812
rect 18966 24760 18972 24812
rect 19024 24760 19030 24812
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19518 24800 19524 24812
rect 19107 24772 19524 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19518 24760 19524 24772
rect 19576 24760 19582 24812
rect 19812 24809 19840 24840
rect 20070 24828 20076 24840
rect 20128 24828 20134 24880
rect 22554 24828 22560 24880
rect 22612 24828 22618 24880
rect 23750 24828 23756 24880
rect 23808 24877 23814 24880
rect 23808 24871 23871 24877
rect 23808 24837 23825 24871
rect 23859 24837 23871 24871
rect 23808 24831 23871 24837
rect 23808 24828 23814 24831
rect 24026 24828 24032 24880
rect 24084 24868 24090 24880
rect 24136 24868 24164 24899
rect 24084 24840 24164 24868
rect 24084 24828 24090 24840
rect 25130 24828 25136 24880
rect 25188 24828 25194 24880
rect 27341 24871 27399 24877
rect 27341 24837 27353 24871
rect 27387 24868 27399 24871
rect 27522 24868 27528 24880
rect 27387 24840 27528 24868
rect 27387 24837 27399 24840
rect 27341 24831 27399 24837
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 19797 24803 19855 24809
rect 19797 24769 19809 24803
rect 19843 24769 19855 24803
rect 19797 24763 19855 24769
rect 19978 24760 19984 24812
rect 20036 24800 20042 24812
rect 21726 24800 21732 24812
rect 20036 24772 21732 24800
rect 20036 24760 20042 24772
rect 21726 24760 21732 24772
rect 21784 24800 21790 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21784 24772 21833 24800
rect 21784 24760 21790 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 23492 24772 23980 24800
rect 22097 24735 22155 24741
rect 12360 24704 20024 24732
rect 7558 24664 7564 24676
rect 5684 24636 6776 24664
rect 6840 24636 7564 24664
rect 5684 24624 5690 24636
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 2406 24596 2412 24608
rect 1627 24568 2412 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 5997 24599 6055 24605
rect 5997 24565 6009 24599
rect 6043 24596 6055 24599
rect 6086 24596 6092 24608
rect 6043 24568 6092 24596
rect 6043 24565 6055 24568
rect 5997 24559 6055 24565
rect 6086 24556 6092 24568
rect 6144 24556 6150 24608
rect 6748 24596 6776 24636
rect 7558 24624 7564 24636
rect 7616 24624 7622 24676
rect 7650 24624 7656 24676
rect 7708 24664 7714 24676
rect 7708 24636 10180 24664
rect 7708 24624 7714 24636
rect 6917 24599 6975 24605
rect 6917 24596 6929 24599
rect 6748 24568 6929 24596
rect 6917 24565 6929 24568
rect 6963 24565 6975 24599
rect 6917 24559 6975 24565
rect 8113 24599 8171 24605
rect 8113 24565 8125 24599
rect 8159 24596 8171 24599
rect 8938 24596 8944 24608
rect 8159 24568 8944 24596
rect 8159 24565 8171 24568
rect 8113 24559 8171 24565
rect 8938 24556 8944 24568
rect 8996 24556 9002 24608
rect 9950 24556 9956 24608
rect 10008 24556 10014 24608
rect 10152 24596 10180 24636
rect 10226 24624 10232 24676
rect 10284 24664 10290 24676
rect 10284 24636 14872 24664
rect 10284 24624 10290 24636
rect 11146 24596 11152 24608
rect 10152 24568 11152 24596
rect 11146 24556 11152 24568
rect 11204 24596 11210 24608
rect 11974 24596 11980 24608
rect 11204 24568 11980 24596
rect 11204 24556 11210 24568
rect 11974 24556 11980 24568
rect 12032 24556 12038 24608
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 14734 24596 14740 24608
rect 14608 24568 14740 24596
rect 14608 24556 14614 24568
rect 14734 24556 14740 24568
rect 14792 24556 14798 24608
rect 14844 24596 14872 24636
rect 15470 24624 15476 24676
rect 15528 24664 15534 24676
rect 16942 24664 16948 24676
rect 15528 24636 16948 24664
rect 15528 24624 15534 24636
rect 16942 24624 16948 24636
rect 17000 24664 17006 24676
rect 17310 24664 17316 24676
rect 17000 24636 17316 24664
rect 17000 24624 17006 24636
rect 17310 24624 17316 24636
rect 17368 24624 17374 24676
rect 17494 24624 17500 24676
rect 17552 24664 17558 24676
rect 19150 24664 19156 24676
rect 17552 24636 19156 24664
rect 17552 24624 17558 24636
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 19702 24624 19708 24676
rect 19760 24664 19766 24676
rect 19889 24667 19947 24673
rect 19889 24664 19901 24667
rect 19760 24636 19901 24664
rect 19760 24624 19766 24636
rect 19889 24633 19901 24636
rect 19935 24633 19947 24667
rect 19889 24627 19947 24633
rect 16574 24596 16580 24608
rect 14844 24568 16580 24596
rect 16574 24556 16580 24568
rect 16632 24556 16638 24608
rect 17129 24599 17187 24605
rect 17129 24565 17141 24599
rect 17175 24596 17187 24599
rect 17586 24596 17592 24608
rect 17175 24568 17592 24596
rect 17175 24565 17187 24568
rect 17129 24559 17187 24565
rect 17586 24556 17592 24568
rect 17644 24556 17650 24608
rect 17678 24556 17684 24608
rect 17736 24556 17742 24608
rect 19245 24599 19303 24605
rect 19245 24565 19257 24599
rect 19291 24596 19303 24599
rect 19610 24596 19616 24608
rect 19291 24568 19616 24596
rect 19291 24565 19303 24568
rect 19245 24559 19303 24565
rect 19610 24556 19616 24568
rect 19668 24556 19674 24608
rect 19996 24596 20024 24704
rect 22097 24701 22109 24735
rect 22143 24732 22155 24735
rect 22830 24732 22836 24744
rect 22143 24704 22836 24732
rect 22143 24701 22155 24704
rect 22097 24695 22155 24701
rect 22830 24692 22836 24704
rect 22888 24692 22894 24744
rect 20070 24624 20076 24676
rect 20128 24664 20134 24676
rect 20622 24664 20628 24676
rect 20128 24636 20628 24664
rect 20128 24624 20134 24636
rect 20622 24624 20628 24636
rect 20680 24664 20686 24676
rect 21818 24664 21824 24676
rect 20680 24636 21824 24664
rect 20680 24624 20686 24636
rect 21818 24624 21824 24636
rect 21876 24624 21882 24676
rect 23492 24596 23520 24772
rect 23566 24692 23572 24744
rect 23624 24692 23630 24744
rect 23584 24664 23612 24692
rect 23952 24664 23980 24772
rect 26234 24760 26240 24812
rect 26292 24760 26298 24812
rect 27154 24760 27160 24812
rect 27212 24800 27218 24812
rect 27249 24803 27307 24809
rect 27249 24800 27261 24803
rect 27212 24772 27261 24800
rect 27212 24760 27218 24772
rect 27249 24769 27261 24772
rect 27295 24769 27307 24803
rect 27249 24763 27307 24769
rect 27430 24760 27436 24812
rect 27488 24760 27494 24812
rect 27614 24760 27620 24812
rect 27672 24760 27678 24812
rect 29270 24760 29276 24812
rect 29328 24760 29334 24812
rect 24210 24692 24216 24744
rect 24268 24732 24274 24744
rect 25593 24735 25651 24741
rect 25593 24732 25605 24735
rect 24268 24704 25605 24732
rect 24268 24692 24274 24704
rect 25593 24701 25605 24704
rect 25639 24701 25651 24735
rect 25593 24695 25651 24701
rect 25869 24735 25927 24741
rect 25869 24701 25881 24735
rect 25915 24732 25927 24735
rect 27632 24732 27660 24760
rect 25915 24704 27660 24732
rect 25915 24701 25927 24704
rect 25869 24695 25927 24701
rect 27617 24667 27675 24673
rect 23584 24636 23888 24664
rect 23952 24636 24256 24664
rect 19996 24568 23520 24596
rect 23658 24556 23664 24608
rect 23716 24556 23722 24608
rect 23860 24605 23888 24636
rect 23845 24599 23903 24605
rect 23845 24565 23857 24599
rect 23891 24565 23903 24599
rect 24228 24596 24256 24636
rect 25792 24636 27200 24664
rect 25792 24596 25820 24636
rect 24228 24568 25820 24596
rect 23845 24559 23903 24565
rect 26326 24556 26332 24608
rect 26384 24556 26390 24608
rect 26786 24556 26792 24608
rect 26844 24596 26850 24608
rect 27065 24599 27123 24605
rect 27065 24596 27077 24599
rect 26844 24568 27077 24596
rect 26844 24556 26850 24568
rect 27065 24565 27077 24568
rect 27111 24565 27123 24599
rect 27172 24596 27200 24636
rect 27617 24633 27629 24667
rect 27663 24664 27675 24667
rect 27798 24664 27804 24676
rect 27663 24636 27804 24664
rect 27663 24633 27675 24636
rect 27617 24627 27675 24633
rect 27798 24624 27804 24636
rect 27856 24624 27862 24676
rect 29181 24599 29239 24605
rect 29181 24596 29193 24599
rect 27172 24568 29193 24596
rect 27065 24559 27123 24565
rect 29181 24565 29193 24568
rect 29227 24565 29239 24599
rect 29181 24559 29239 24565
rect 1104 24506 29716 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 29716 24506
rect 1104 24432 29716 24454
rect 2120 24395 2178 24401
rect 2120 24361 2132 24395
rect 2166 24392 2178 24395
rect 3973 24395 4031 24401
rect 3973 24392 3985 24395
rect 2166 24364 3985 24392
rect 2166 24361 2178 24364
rect 2120 24355 2178 24361
rect 3973 24361 3985 24364
rect 4019 24361 4031 24395
rect 3973 24355 4031 24361
rect 4157 24395 4215 24401
rect 4157 24361 4169 24395
rect 4203 24392 4215 24395
rect 4985 24395 5043 24401
rect 4985 24392 4997 24395
rect 4203 24364 4997 24392
rect 4203 24361 4215 24364
rect 4157 24355 4215 24361
rect 4985 24361 4997 24364
rect 5031 24361 5043 24395
rect 4985 24355 5043 24361
rect 5350 24352 5356 24404
rect 5408 24352 5414 24404
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 6270 24392 6276 24404
rect 5592 24364 6276 24392
rect 5592 24352 5598 24364
rect 6270 24352 6276 24364
rect 6328 24352 6334 24404
rect 7558 24352 7564 24404
rect 7616 24352 7622 24404
rect 7834 24392 7840 24404
rect 7668 24364 7840 24392
rect 4246 24284 4252 24336
rect 4304 24324 4310 24336
rect 4525 24327 4583 24333
rect 4525 24324 4537 24327
rect 4304 24296 4537 24324
rect 4304 24284 4310 24296
rect 4525 24293 4537 24296
rect 4571 24324 4583 24327
rect 4798 24324 4804 24336
rect 4571 24296 4804 24324
rect 4571 24293 4583 24296
rect 4525 24287 4583 24293
rect 4798 24284 4804 24296
rect 4856 24284 4862 24336
rect 5166 24284 5172 24336
rect 5224 24324 5230 24336
rect 5224 24296 6316 24324
rect 5224 24284 5230 24296
rect 1857 24259 1915 24265
rect 1857 24225 1869 24259
rect 1903 24256 1915 24259
rect 2774 24256 2780 24268
rect 1903 24228 2780 24256
rect 1903 24225 1915 24228
rect 1857 24219 1915 24225
rect 2774 24216 2780 24228
rect 2832 24256 2838 24268
rect 3694 24256 3700 24268
rect 2832 24228 3700 24256
rect 2832 24216 2838 24228
rect 3694 24216 3700 24228
rect 3752 24216 3758 24268
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 4614 24256 4620 24268
rect 4212 24228 4620 24256
rect 4212 24216 4218 24228
rect 4614 24216 4620 24228
rect 4672 24256 4678 24268
rect 4672 24228 4936 24256
rect 4672 24216 4678 24228
rect 3234 24148 3240 24200
rect 3292 24148 3298 24200
rect 4522 24148 4528 24200
rect 4580 24188 4586 24200
rect 4908 24197 4936 24228
rect 5092 24228 5488 24256
rect 5092 24197 5120 24228
rect 5460 24197 5488 24228
rect 6178 24216 6184 24268
rect 6236 24216 6242 24268
rect 4801 24191 4859 24197
rect 4801 24188 4813 24191
rect 4580 24160 4813 24188
rect 4580 24148 4586 24160
rect 4801 24157 4813 24160
rect 4847 24157 4859 24191
rect 4801 24151 4859 24157
rect 4893 24191 4951 24197
rect 4893 24157 4905 24191
rect 4939 24157 4951 24191
rect 4893 24151 4951 24157
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5077 24151 5135 24157
rect 5261 24191 5319 24197
rect 5261 24157 5273 24191
rect 5307 24157 5319 24191
rect 5261 24151 5319 24157
rect 5445 24191 5503 24197
rect 5445 24157 5457 24191
rect 5491 24188 5503 24191
rect 5534 24188 5540 24200
rect 5491 24160 5540 24188
rect 5491 24157 5503 24160
rect 5445 24151 5503 24157
rect 4540 24120 4568 24148
rect 3620 24092 4568 24120
rect 4709 24123 4767 24129
rect 3620 24061 3648 24092
rect 4709 24089 4721 24123
rect 4755 24120 4767 24123
rect 5092 24120 5120 24151
rect 4755 24092 5120 24120
rect 5276 24120 5304 24151
rect 5534 24148 5540 24160
rect 5592 24148 5598 24200
rect 5902 24148 5908 24200
rect 5960 24148 5966 24200
rect 6053 24191 6111 24197
rect 6053 24157 6065 24191
rect 6099 24188 6111 24191
rect 6196 24188 6224 24216
rect 6288 24197 6316 24296
rect 6730 24284 6736 24336
rect 6788 24324 6794 24336
rect 7668 24324 7696 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 8202 24352 8208 24404
rect 8260 24392 8266 24404
rect 9950 24392 9956 24404
rect 8260 24364 9956 24392
rect 8260 24352 8266 24364
rect 6788 24296 7696 24324
rect 7760 24296 8432 24324
rect 6788 24284 6794 24296
rect 7760 24200 7788 24296
rect 8202 24256 8208 24268
rect 7852 24228 8208 24256
rect 6099 24160 6224 24188
rect 6273 24191 6331 24197
rect 6099 24157 6111 24160
rect 6053 24151 6111 24157
rect 6273 24157 6285 24191
rect 6319 24157 6331 24191
rect 6273 24151 6331 24157
rect 6370 24191 6428 24197
rect 6370 24157 6382 24191
rect 6416 24157 6428 24191
rect 6370 24151 6428 24157
rect 6178 24120 6184 24132
rect 5276 24092 6184 24120
rect 4755 24089 4767 24092
rect 4709 24083 4767 24089
rect 3605 24055 3663 24061
rect 3605 24021 3617 24055
rect 3651 24021 3663 24055
rect 3605 24015 3663 24021
rect 3878 24012 3884 24064
rect 3936 24052 3942 24064
rect 4157 24055 4215 24061
rect 4157 24052 4169 24055
rect 3936 24024 4169 24052
rect 3936 24012 3942 24024
rect 4157 24021 4169 24024
rect 4203 24021 4215 24055
rect 4157 24015 4215 24021
rect 4338 24012 4344 24064
rect 4396 24052 4402 24064
rect 4724 24052 4752 24083
rect 6178 24080 6184 24092
rect 6236 24080 6242 24132
rect 4396 24024 4752 24052
rect 4396 24012 4402 24024
rect 5994 24012 6000 24064
rect 6052 24052 6058 24064
rect 6380 24052 6408 24151
rect 7742 24148 7748 24200
rect 7800 24148 7806 24200
rect 7852 24197 7880 24228
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 7837 24191 7895 24197
rect 7837 24157 7849 24191
rect 7883 24157 7895 24191
rect 7837 24151 7895 24157
rect 8110 24148 8116 24200
rect 8168 24148 8174 24200
rect 8404 24197 8432 24296
rect 8588 24197 8616 24364
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 13906 24352 13912 24404
rect 13964 24392 13970 24404
rect 13964 24364 14872 24392
rect 13964 24352 13970 24364
rect 8665 24327 8723 24333
rect 8665 24293 8677 24327
rect 8711 24324 8723 24327
rect 8754 24324 8760 24336
rect 8711 24296 8760 24324
rect 8711 24293 8723 24296
rect 8665 24287 8723 24293
rect 8754 24284 8760 24296
rect 8812 24284 8818 24336
rect 9585 24327 9643 24333
rect 9585 24293 9597 24327
rect 9631 24324 9643 24327
rect 14458 24324 14464 24336
rect 9631 24296 14464 24324
rect 9631 24293 9643 24296
rect 9585 24287 9643 24293
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 14737 24327 14795 24333
rect 14737 24293 14749 24327
rect 14783 24293 14795 24327
rect 14844 24324 14872 24364
rect 14918 24352 14924 24404
rect 14976 24392 14982 24404
rect 16850 24392 16856 24404
rect 14976 24364 16856 24392
rect 14976 24352 14982 24364
rect 16850 24352 16856 24364
rect 16908 24352 16914 24404
rect 16942 24352 16948 24404
rect 17000 24392 17006 24404
rect 17402 24392 17408 24404
rect 17000 24364 17408 24392
rect 17000 24352 17006 24364
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 17586 24352 17592 24404
rect 17644 24392 17650 24404
rect 18230 24392 18236 24404
rect 17644 24364 18236 24392
rect 17644 24352 17650 24364
rect 18230 24352 18236 24364
rect 18288 24392 18294 24404
rect 18288 24364 19288 24392
rect 18288 24352 18294 24364
rect 15010 24324 15016 24336
rect 14844 24296 15016 24324
rect 14737 24287 14795 24293
rect 8846 24216 8852 24268
rect 8904 24256 8910 24268
rect 10226 24256 10232 24268
rect 8904 24228 9352 24256
rect 8904 24216 8910 24228
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 8541 24191 8616 24197
rect 8541 24157 8553 24191
rect 8587 24160 8616 24191
rect 8587 24157 8599 24160
rect 8541 24151 8599 24157
rect 8662 24148 8668 24200
rect 8720 24188 8726 24200
rect 8757 24191 8815 24197
rect 8757 24188 8769 24191
rect 8720 24160 8769 24188
rect 8720 24148 8726 24160
rect 8757 24157 8769 24160
rect 8803 24157 8815 24191
rect 8757 24151 8815 24157
rect 8938 24148 8944 24200
rect 8996 24148 9002 24200
rect 9324 24197 9352 24228
rect 9876 24228 10232 24256
rect 9125 24191 9183 24197
rect 9125 24157 9137 24191
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9217 24151 9275 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 9677 24191 9735 24197
rect 9677 24157 9689 24191
rect 9723 24188 9735 24191
rect 9766 24188 9772 24200
rect 9723 24160 9772 24188
rect 9723 24157 9735 24160
rect 9677 24151 9735 24157
rect 7926 24080 7932 24132
rect 7984 24080 7990 24132
rect 8205 24123 8263 24129
rect 8205 24089 8217 24123
rect 8251 24120 8263 24123
rect 9140 24120 9168 24151
rect 8251 24092 9168 24120
rect 8251 24089 8263 24092
rect 8205 24083 8263 24089
rect 6052 24024 6408 24052
rect 6549 24055 6607 24061
rect 6052 24012 6058 24024
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 9232 24052 9260 24151
rect 9766 24148 9772 24160
rect 9824 24148 9830 24200
rect 9876 24197 9904 24228
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 10410 24256 10416 24268
rect 10336 24228 10416 24256
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 9950 24148 9956 24200
rect 10008 24148 10014 24200
rect 10336 24197 10364 24228
rect 10410 24216 10416 24228
rect 10468 24216 10474 24268
rect 11900 24228 12664 24256
rect 11900 24197 11928 24228
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24157 10379 24191
rect 10689 24191 10747 24197
rect 10689 24188 10701 24191
rect 10321 24151 10379 24157
rect 10428 24160 10701 24188
rect 10060 24120 10088 24151
rect 10428 24120 10456 24160
rect 10689 24157 10701 24160
rect 10735 24157 10747 24191
rect 10689 24151 10747 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 11974 24148 11980 24200
rect 12032 24188 12038 24200
rect 12032 24160 12077 24188
rect 12032 24148 12038 24160
rect 12158 24148 12164 24200
rect 12216 24148 12222 24200
rect 12250 24148 12256 24200
rect 12308 24148 12314 24200
rect 12350 24191 12408 24197
rect 12350 24157 12362 24191
rect 12396 24188 12408 24191
rect 12526 24188 12532 24200
rect 12396 24160 12532 24188
rect 12396 24157 12408 24160
rect 12350 24151 12408 24157
rect 9968 24092 10088 24120
rect 10152 24092 10456 24120
rect 9968 24064 9996 24092
rect 6595 24024 9260 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 9950 24012 9956 24064
rect 10008 24012 10014 24064
rect 10042 24012 10048 24064
rect 10100 24052 10106 24064
rect 10152 24052 10180 24092
rect 10502 24080 10508 24132
rect 10560 24080 10566 24132
rect 10594 24080 10600 24132
rect 10652 24080 10658 24132
rect 11606 24080 11612 24132
rect 11664 24120 11670 24132
rect 12360 24120 12388 24151
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 11664 24092 12388 24120
rect 11664 24080 11670 24092
rect 10100 24024 10180 24052
rect 10100 24012 10106 24024
rect 10226 24012 10232 24064
rect 10284 24012 10290 24064
rect 10778 24012 10784 24064
rect 10836 24052 10842 24064
rect 10873 24055 10931 24061
rect 10873 24052 10885 24055
rect 10836 24024 10885 24052
rect 10836 24012 10842 24024
rect 10873 24021 10885 24024
rect 10919 24021 10931 24055
rect 10873 24015 10931 24021
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 12636 24061 12664 24228
rect 13906 24216 13912 24268
rect 13964 24256 13970 24268
rect 14090 24256 14096 24268
rect 13964 24228 14096 24256
rect 13964 24216 13970 24228
rect 14090 24216 14096 24228
rect 14148 24216 14154 24268
rect 14185 24259 14243 24265
rect 14185 24225 14197 24259
rect 14231 24256 14243 24259
rect 14752 24256 14780 24287
rect 15010 24284 15016 24296
rect 15068 24284 15074 24336
rect 15749 24327 15807 24333
rect 15749 24293 15761 24327
rect 15795 24324 15807 24327
rect 18414 24324 18420 24336
rect 15795 24296 18420 24324
rect 15795 24293 15807 24296
rect 15749 24287 15807 24293
rect 18414 24284 18420 24296
rect 18472 24284 18478 24336
rect 19260 24324 19288 24364
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 22465 24395 22523 24401
rect 19392 24364 21772 24392
rect 19392 24352 19398 24364
rect 19978 24324 19984 24336
rect 19260 24296 19984 24324
rect 18785 24259 18843 24265
rect 14231 24228 14688 24256
rect 14752 24228 18644 24256
rect 14231 24225 14243 24228
rect 14185 24219 14243 24225
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24188 12863 24191
rect 13173 24191 13231 24197
rect 12851 24160 13124 24188
rect 12851 24157 12863 24160
rect 12805 24151 12863 24157
rect 12894 24080 12900 24132
rect 12952 24080 12958 24132
rect 12986 24080 12992 24132
rect 13044 24080 13050 24132
rect 13096 24120 13124 24160
rect 13173 24157 13185 24191
rect 13219 24188 13231 24191
rect 13262 24188 13268 24200
rect 13219 24160 13268 24188
rect 13219 24157 13231 24160
rect 13173 24151 13231 24157
rect 13262 24148 13268 24160
rect 13320 24148 13326 24200
rect 14556 24191 14614 24197
rect 14556 24188 14568 24191
rect 14292 24160 14568 24188
rect 13538 24120 13544 24132
rect 13096 24092 13544 24120
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 13998 24080 14004 24132
rect 14056 24120 14062 24132
rect 14292 24120 14320 24160
rect 14556 24157 14568 24160
rect 14602 24157 14614 24191
rect 14660 24188 14688 24228
rect 14660 24160 14872 24188
rect 14556 24151 14614 24157
rect 14844 24132 14872 24160
rect 15010 24148 15016 24200
rect 15068 24148 15074 24200
rect 15286 24148 15292 24200
rect 15344 24148 15350 24200
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15562 24188 15568 24200
rect 15427 24160 15568 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 15654 24148 15660 24200
rect 15712 24148 15718 24200
rect 15838 24148 15844 24200
rect 15896 24148 15902 24200
rect 16850 24148 16856 24200
rect 16908 24148 16914 24200
rect 16942 24148 16948 24200
rect 17000 24148 17006 24200
rect 17218 24197 17224 24200
rect 17201 24191 17224 24197
rect 17201 24157 17213 24191
rect 17276 24190 17282 24200
rect 17276 24162 17356 24190
rect 17201 24151 17224 24157
rect 17218 24148 17224 24151
rect 17276 24148 17282 24162
rect 14056 24092 14320 24120
rect 14056 24080 14062 24092
rect 14826 24080 14832 24132
rect 14884 24120 14890 24132
rect 15197 24123 15255 24129
rect 15197 24120 15209 24123
rect 14884 24092 15209 24120
rect 14884 24080 14890 24092
rect 15197 24089 15209 24092
rect 15243 24089 15255 24123
rect 15197 24083 15255 24089
rect 15580 24092 16988 24120
rect 12529 24055 12587 24061
rect 12529 24052 12541 24055
rect 12492 24024 12541 24052
rect 12492 24012 12498 24024
rect 12529 24021 12541 24024
rect 12575 24021 12587 24055
rect 12529 24015 12587 24021
rect 12621 24055 12679 24061
rect 12621 24021 12633 24055
rect 12667 24052 12679 24055
rect 13078 24052 13084 24064
rect 12667 24024 13084 24052
rect 12667 24021 12679 24024
rect 12621 24015 12679 24021
rect 13078 24012 13084 24024
rect 13136 24012 13142 24064
rect 13262 24012 13268 24064
rect 13320 24052 13326 24064
rect 13722 24052 13728 24064
rect 13320 24024 13728 24052
rect 13320 24012 13326 24024
rect 13722 24012 13728 24024
rect 13780 24052 13786 24064
rect 15580 24061 15608 24092
rect 16960 24064 16988 24092
rect 17034 24080 17040 24132
rect 17092 24080 17098 24132
rect 17328 24120 17356 24162
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 17497 24191 17555 24197
rect 17497 24188 17509 24191
rect 17460 24160 17509 24188
rect 17460 24148 17466 24160
rect 17497 24157 17509 24160
rect 17543 24188 17555 24191
rect 17586 24188 17592 24200
rect 17543 24160 17592 24188
rect 17543 24157 17555 24160
rect 17497 24151 17555 24157
rect 17586 24148 17592 24160
rect 17644 24148 17650 24200
rect 18046 24148 18052 24200
rect 18104 24148 18110 24200
rect 18414 24148 18420 24200
rect 18472 24148 18478 24200
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 18616 24188 18644 24228
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 19334 24256 19340 24268
rect 18831 24228 19340 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 19334 24216 19340 24228
rect 19392 24216 19398 24268
rect 18555 24160 18644 24188
rect 18877 24191 18935 24197
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 18877 24157 18889 24191
rect 18923 24157 18935 24191
rect 19444 24188 19472 24296
rect 19978 24284 19984 24296
rect 20036 24284 20042 24336
rect 21082 24324 21088 24336
rect 20088 24296 21088 24324
rect 19797 24259 19855 24265
rect 19797 24225 19809 24259
rect 19843 24256 19855 24259
rect 20088 24256 20116 24296
rect 21082 24284 21088 24296
rect 21140 24284 21146 24336
rect 19843 24228 20116 24256
rect 20441 24259 20499 24265
rect 19843 24225 19855 24228
rect 19797 24219 19855 24225
rect 20441 24225 20453 24259
rect 20487 24256 20499 24259
rect 21637 24259 21695 24265
rect 21637 24256 21649 24259
rect 20487 24228 21649 24256
rect 20487 24225 20499 24228
rect 20441 24219 20499 24225
rect 21637 24225 21649 24228
rect 21683 24225 21695 24259
rect 21637 24219 21695 24225
rect 19613 24191 19671 24197
rect 19613 24188 19625 24191
rect 19444 24160 19625 24188
rect 18877 24151 18935 24157
rect 19613 24157 19625 24160
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 17957 24123 18015 24129
rect 17957 24120 17969 24123
rect 17328 24092 17969 24120
rect 17957 24089 17969 24092
rect 18003 24120 18015 24123
rect 18892 24120 18920 24151
rect 19702 24148 19708 24200
rect 19760 24188 19766 24200
rect 19889 24191 19947 24197
rect 19889 24188 19901 24191
rect 19760 24160 19901 24188
rect 19760 24148 19766 24160
rect 19889 24157 19901 24160
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24188 20223 24191
rect 20456 24188 20484 24219
rect 20533 24194 20591 24197
rect 20211 24160 20484 24188
rect 20211 24157 20223 24160
rect 20165 24151 20223 24157
rect 18003 24092 18920 24120
rect 18003 24089 18015 24092
rect 17957 24083 18015 24089
rect 19242 24080 19248 24132
rect 19300 24120 19306 24132
rect 19996 24120 20024 24151
rect 20530 24142 20536 24194
rect 20588 24142 20594 24194
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20732 24160 21005 24188
rect 19300 24092 20024 24120
rect 19300 24080 19306 24092
rect 20070 24080 20076 24132
rect 20128 24120 20134 24132
rect 20128 24092 20484 24120
rect 20128 24080 20134 24092
rect 14553 24055 14611 24061
rect 14553 24052 14565 24055
rect 13780 24024 14565 24052
rect 13780 24012 13786 24024
rect 14553 24021 14565 24024
rect 14599 24021 14611 24055
rect 14553 24015 14611 24021
rect 15565 24055 15623 24061
rect 15565 24021 15577 24055
rect 15611 24021 15623 24055
rect 15565 24015 15623 24021
rect 16666 24012 16672 24064
rect 16724 24012 16730 24064
rect 16942 24012 16948 24064
rect 17000 24012 17006 24064
rect 18138 24012 18144 24064
rect 18196 24012 18202 24064
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 18647 24024 19441 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 19429 24021 19441 24024
rect 19475 24052 19487 24055
rect 19702 24052 19708 24064
rect 19475 24024 19708 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 19702 24012 19708 24024
rect 19760 24012 19766 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 20257 24055 20315 24061
rect 20257 24052 20269 24055
rect 19944 24024 20269 24052
rect 19944 24012 19950 24024
rect 20257 24021 20269 24024
rect 20303 24021 20315 24055
rect 20456 24052 20484 24092
rect 20732 24052 20760 24160
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 20993 24151 21051 24157
rect 21358 24148 21364 24200
rect 21416 24148 21422 24200
rect 21082 24080 21088 24132
rect 21140 24120 21146 24132
rect 21177 24123 21235 24129
rect 21177 24120 21189 24123
rect 21140 24092 21189 24120
rect 21140 24080 21146 24092
rect 21177 24089 21189 24092
rect 21223 24089 21235 24123
rect 21177 24083 21235 24089
rect 21266 24080 21272 24132
rect 21324 24120 21330 24132
rect 21744 24120 21772 24364
rect 22465 24361 22477 24395
rect 22511 24392 22523 24395
rect 22554 24392 22560 24404
rect 22511 24364 22560 24392
rect 22511 24361 22523 24364
rect 22465 24355 22523 24361
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 22925 24395 22983 24401
rect 22925 24392 22937 24395
rect 22888 24364 22937 24392
rect 22888 24352 22894 24364
rect 22925 24361 22937 24364
rect 22971 24361 22983 24395
rect 22925 24355 22983 24361
rect 24210 24352 24216 24404
rect 24268 24352 24274 24404
rect 25130 24352 25136 24404
rect 25188 24392 25194 24404
rect 25225 24395 25283 24401
rect 25225 24392 25237 24395
rect 25188 24364 25237 24392
rect 25188 24352 25194 24364
rect 25225 24361 25237 24364
rect 25271 24361 25283 24395
rect 26234 24392 26240 24404
rect 25225 24355 25283 24361
rect 25424 24364 26240 24392
rect 21818 24284 21824 24336
rect 21876 24284 21882 24336
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 22060 24296 22416 24324
rect 22060 24284 22066 24296
rect 21836 24256 21864 24284
rect 21836 24228 22048 24256
rect 21818 24148 21824 24200
rect 21876 24148 21882 24200
rect 21910 24148 21916 24200
rect 21968 24148 21974 24200
rect 22020 24188 22048 24228
rect 22094 24216 22100 24268
rect 22152 24216 22158 24268
rect 22388 24197 22416 24296
rect 23106 24284 23112 24336
rect 23164 24284 23170 24336
rect 25424 24324 25452 24364
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 27157 24395 27215 24401
rect 27157 24361 27169 24395
rect 27203 24392 27215 24395
rect 27430 24392 27436 24404
rect 27203 24364 27436 24392
rect 27203 24361 27215 24364
rect 27157 24355 27215 24361
rect 27430 24352 27436 24364
rect 27488 24352 27494 24404
rect 23676 24296 25452 24324
rect 22189 24191 22247 24197
rect 22189 24188 22201 24191
rect 22020 24160 22201 24188
rect 22189 24157 22201 24160
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 22373 24191 22431 24197
rect 22373 24157 22385 24191
rect 22419 24188 22431 24191
rect 23676 24188 23704 24296
rect 23750 24216 23756 24268
rect 23808 24216 23814 24268
rect 22419 24160 23704 24188
rect 23845 24191 23903 24197
rect 22419 24157 22431 24160
rect 22373 24151 22431 24157
rect 23845 24157 23857 24191
rect 23891 24188 23903 24191
rect 24026 24188 24032 24200
rect 23891 24160 24032 24188
rect 23891 24157 23903 24160
rect 23845 24151 23903 24157
rect 24026 24148 24032 24160
rect 24084 24148 24090 24200
rect 25332 24197 25360 24296
rect 25409 24259 25467 24265
rect 25409 24225 25421 24259
rect 25455 24256 25467 24259
rect 25455 24228 27660 24256
rect 25455 24225 25467 24228
rect 25409 24219 25467 24225
rect 27632 24200 27660 24228
rect 25317 24191 25375 24197
rect 25317 24157 25329 24191
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 27614 24148 27620 24200
rect 27672 24148 27678 24200
rect 23385 24123 23443 24129
rect 21324 24092 21680 24120
rect 21744 24092 22094 24120
rect 21324 24080 21330 24092
rect 20456 24024 20760 24052
rect 20257 24015 20315 24021
rect 20898 24012 20904 24064
rect 20956 24012 20962 24064
rect 21542 24012 21548 24064
rect 21600 24012 21606 24064
rect 21652 24052 21680 24092
rect 21910 24052 21916 24064
rect 21652 24024 21916 24052
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 22066 24052 22094 24092
rect 23385 24089 23397 24123
rect 23431 24120 23443 24123
rect 23658 24120 23664 24132
rect 23431 24092 23664 24120
rect 23431 24089 23443 24092
rect 23385 24083 23443 24089
rect 23658 24080 23664 24092
rect 23716 24120 23722 24132
rect 23934 24120 23940 24132
rect 23716 24092 23940 24120
rect 23716 24080 23722 24092
rect 23934 24080 23940 24092
rect 23992 24080 23998 24132
rect 25682 24080 25688 24132
rect 25740 24080 25746 24132
rect 26326 24080 26332 24132
rect 26384 24080 26390 24132
rect 27893 24123 27951 24129
rect 27893 24089 27905 24123
rect 27939 24120 27951 24123
rect 28166 24120 28172 24132
rect 27939 24092 28172 24120
rect 27939 24089 27951 24092
rect 27893 24083 27951 24089
rect 28166 24080 28172 24092
rect 28224 24080 28230 24132
rect 28902 24080 28908 24132
rect 28960 24080 28966 24132
rect 26510 24052 26516 24064
rect 22066 24024 26516 24052
rect 26510 24012 26516 24024
rect 26568 24012 26574 24064
rect 27522 24012 27528 24064
rect 27580 24052 27586 24064
rect 29365 24055 29423 24061
rect 29365 24052 29377 24055
rect 27580 24024 29377 24052
rect 27580 24012 27586 24024
rect 29365 24021 29377 24024
rect 29411 24021 29423 24055
rect 29365 24015 29423 24021
rect 1104 23962 29716 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 29716 23962
rect 1104 23888 29716 23910
rect 3234 23808 3240 23860
rect 3292 23808 3298 23860
rect 4246 23808 4252 23860
rect 4304 23808 4310 23860
rect 4617 23851 4675 23857
rect 4617 23817 4629 23851
rect 4663 23848 4675 23851
rect 4798 23848 4804 23860
rect 4663 23820 4804 23848
rect 4663 23817 4675 23820
rect 4617 23811 4675 23817
rect 4798 23808 4804 23820
rect 4856 23808 4862 23860
rect 7650 23808 7656 23860
rect 7708 23848 7714 23860
rect 7745 23851 7803 23857
rect 7745 23848 7757 23851
rect 7708 23820 7757 23848
rect 7708 23808 7714 23820
rect 7745 23817 7757 23820
rect 7791 23817 7803 23851
rect 7745 23811 7803 23817
rect 8018 23808 8024 23860
rect 8076 23848 8082 23860
rect 9861 23851 9919 23857
rect 8076 23820 8800 23848
rect 8076 23808 8082 23820
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 4985 23783 5043 23789
rect 4580 23752 4844 23780
rect 4580 23740 4586 23752
rect 842 23672 848 23724
rect 900 23712 906 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 900 23684 1409 23712
rect 900 23672 906 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23712 3387 23715
rect 3970 23712 3976 23724
rect 3375 23684 3976 23712
rect 3375 23681 3387 23684
rect 3329 23675 3387 23681
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 4154 23672 4160 23724
rect 4212 23672 4218 23724
rect 4338 23672 4344 23724
rect 4396 23672 4402 23724
rect 4816 23721 4844 23752
rect 4985 23749 4997 23783
rect 5031 23780 5043 23783
rect 5258 23780 5264 23792
rect 5031 23752 5264 23780
rect 5031 23749 5043 23752
rect 4985 23743 5043 23749
rect 5258 23740 5264 23752
rect 5316 23780 5322 23792
rect 5316 23752 7052 23780
rect 5316 23740 5322 23752
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23681 4767 23715
rect 4709 23675 4767 23681
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23712 4859 23715
rect 4890 23712 4896 23724
rect 4847 23684 4896 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 4724 23644 4752 23675
rect 4890 23672 4896 23684
rect 4948 23672 4954 23724
rect 5905 23715 5963 23721
rect 5905 23681 5917 23715
rect 5951 23712 5963 23715
rect 6086 23712 6092 23724
rect 5951 23684 6092 23712
rect 5951 23681 5963 23684
rect 5905 23675 5963 23681
rect 6086 23672 6092 23684
rect 6144 23672 6150 23724
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6546 23712 6552 23724
rect 6328 23684 6552 23712
rect 6328 23672 6334 23684
rect 6546 23672 6552 23684
rect 6604 23712 6610 23724
rect 7024 23721 7052 23752
rect 7392 23752 8708 23780
rect 6641 23715 6699 23721
rect 6641 23712 6653 23715
rect 6604 23684 6653 23712
rect 6604 23672 6610 23684
rect 6641 23681 6653 23684
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 7009 23715 7067 23721
rect 7009 23681 7021 23715
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7190 23672 7196 23724
rect 7248 23672 7254 23724
rect 7392 23721 7420 23752
rect 8680 23724 8708 23752
rect 7285 23715 7343 23721
rect 7285 23681 7297 23715
rect 7331 23681 7343 23715
rect 7285 23675 7343 23681
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 5350 23644 5356 23656
rect 1719 23616 2774 23644
rect 4724 23616 5356 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 2746 23576 2774 23616
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 6362 23604 6368 23656
rect 6420 23644 6426 23656
rect 7300 23644 7328 23675
rect 7558 23672 7564 23724
rect 7616 23712 7622 23724
rect 7653 23715 7711 23721
rect 7653 23712 7665 23715
rect 7616 23684 7665 23712
rect 7616 23672 7622 23684
rect 7653 23681 7665 23684
rect 7699 23681 7711 23715
rect 7653 23675 7711 23681
rect 8018 23672 8024 23724
rect 8076 23712 8082 23724
rect 8297 23715 8355 23721
rect 8297 23712 8309 23715
rect 8076 23684 8309 23712
rect 8076 23672 8082 23684
rect 8297 23681 8309 23684
rect 8343 23681 8355 23715
rect 8570 23712 8576 23724
rect 8297 23675 8355 23681
rect 8404 23684 8576 23712
rect 8404 23644 8432 23684
rect 8570 23672 8576 23684
rect 8628 23672 8634 23724
rect 8662 23672 8668 23724
rect 8720 23672 8726 23724
rect 8772 23712 8800 23820
rect 9861 23817 9873 23851
rect 9907 23848 9919 23851
rect 11333 23851 11391 23857
rect 9907 23820 10272 23848
rect 9907 23817 9919 23820
rect 9861 23811 9919 23817
rect 8849 23783 8907 23789
rect 8849 23749 8861 23783
rect 8895 23780 8907 23783
rect 8895 23752 9812 23780
rect 8895 23749 8907 23752
rect 8849 23743 8907 23749
rect 9784 23724 9812 23752
rect 9309 23715 9367 23721
rect 9309 23712 9321 23715
rect 8772 23684 9321 23712
rect 9309 23681 9321 23684
rect 9355 23681 9367 23715
rect 9309 23675 9367 23681
rect 9398 23672 9404 23724
rect 9456 23712 9462 23724
rect 9493 23715 9551 23721
rect 9493 23712 9505 23715
rect 9456 23684 9505 23712
rect 9456 23672 9462 23684
rect 9493 23681 9505 23684
rect 9539 23681 9551 23715
rect 9493 23675 9551 23681
rect 9582 23672 9588 23724
rect 9640 23672 9646 23724
rect 9674 23672 9680 23724
rect 9732 23672 9738 23724
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 10244 23721 10272 23820
rect 11333 23817 11345 23851
rect 11379 23817 11391 23851
rect 11333 23811 11391 23817
rect 13265 23851 13323 23857
rect 13265 23817 13277 23851
rect 13311 23848 13323 23851
rect 14461 23851 14519 23857
rect 13311 23820 14136 23848
rect 13311 23817 13323 23820
rect 13265 23811 13323 23817
rect 11146 23740 11152 23792
rect 11204 23740 11210 23792
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 9824 23684 9965 23712
rect 9824 23672 9830 23684
rect 9953 23681 9965 23684
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23681 10103 23715
rect 10045 23675 10103 23681
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23712 10287 23715
rect 10505 23715 10563 23721
rect 10505 23712 10517 23715
rect 10275 23684 10517 23712
rect 10275 23681 10287 23684
rect 10229 23675 10287 23681
rect 10505 23681 10517 23684
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 10689 23715 10747 23721
rect 10689 23681 10701 23715
rect 10735 23712 10747 23715
rect 10778 23712 10784 23724
rect 10735 23684 10784 23712
rect 10735 23681 10747 23684
rect 10689 23675 10747 23681
rect 9416 23644 9444 23672
rect 6420 23616 8432 23644
rect 8496 23616 9444 23644
rect 6420 23604 6426 23616
rect 2746 23548 7328 23576
rect 4433 23511 4491 23517
rect 4433 23477 4445 23511
rect 4479 23508 4491 23511
rect 4706 23508 4712 23520
rect 4479 23480 4712 23508
rect 4479 23477 4491 23480
rect 4433 23471 4491 23477
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 5994 23468 6000 23520
rect 6052 23468 6058 23520
rect 6733 23511 6791 23517
rect 6733 23477 6745 23511
rect 6779 23508 6791 23511
rect 6822 23508 6828 23520
rect 6779 23480 6828 23508
rect 6779 23477 6791 23480
rect 6733 23471 6791 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7300 23508 7328 23548
rect 7374 23536 7380 23588
rect 7432 23576 7438 23588
rect 7561 23579 7619 23585
rect 7561 23576 7573 23579
rect 7432 23548 7573 23576
rect 7432 23536 7438 23548
rect 7561 23545 7573 23548
rect 7607 23576 7619 23579
rect 8294 23576 8300 23588
rect 7607 23548 8300 23576
rect 7607 23545 7619 23548
rect 7561 23539 7619 23545
rect 8294 23536 8300 23548
rect 8352 23536 8358 23588
rect 8389 23579 8447 23585
rect 8389 23545 8401 23579
rect 8435 23576 8447 23579
rect 8496 23576 8524 23616
rect 8435 23548 8524 23576
rect 8435 23545 8447 23548
rect 8389 23539 8447 23545
rect 8570 23536 8576 23588
rect 8628 23576 8634 23588
rect 10060 23576 10088 23675
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 11348 23712 11376 23811
rect 12526 23740 12532 23792
rect 12584 23780 12590 23792
rect 14108 23789 14136 23820
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 17954 23848 17960 23860
rect 14507 23820 17960 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 19242 23808 19248 23860
rect 19300 23848 19306 23860
rect 19518 23848 19524 23860
rect 19300 23820 19524 23848
rect 19300 23808 19306 23820
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 19702 23808 19708 23860
rect 19760 23808 19766 23860
rect 25682 23808 25688 23860
rect 25740 23848 25746 23860
rect 26329 23851 26387 23857
rect 26329 23848 26341 23851
rect 25740 23820 26341 23848
rect 25740 23808 25746 23820
rect 26329 23817 26341 23820
rect 26375 23817 26387 23851
rect 26329 23811 26387 23817
rect 28166 23808 28172 23860
rect 28224 23808 28230 23860
rect 28902 23808 28908 23860
rect 28960 23808 28966 23860
rect 12713 23783 12771 23789
rect 12713 23780 12725 23783
rect 12584 23752 12725 23780
rect 12584 23740 12590 23752
rect 12713 23749 12725 23752
rect 12759 23780 12771 23783
rect 14093 23783 14151 23789
rect 12759 23752 13400 23780
rect 12759 23749 12771 23752
rect 12713 23743 12771 23749
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 11348 23684 11529 23712
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23681 11759 23715
rect 11701 23675 11759 23681
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23681 12035 23715
rect 11977 23675 12035 23681
rect 12161 23715 12219 23721
rect 12161 23681 12173 23715
rect 12207 23712 12219 23715
rect 12989 23715 13047 23721
rect 12989 23712 13001 23715
rect 12207 23684 13001 23712
rect 12207 23681 12219 23684
rect 12161 23675 12219 23681
rect 12989 23681 13001 23684
rect 13035 23681 13047 23715
rect 12989 23675 13047 23681
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23644 10471 23647
rect 11716 23644 11744 23675
rect 10459 23616 11744 23644
rect 10459 23613 10471 23616
rect 10413 23607 10471 23613
rect 8628 23548 10088 23576
rect 8628 23536 8634 23548
rect 10226 23536 10232 23588
rect 10284 23576 10290 23588
rect 11992 23576 12020 23675
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 13372 23721 13400 23752
rect 14093 23749 14105 23783
rect 14139 23749 14151 23783
rect 14093 23743 14151 23749
rect 14182 23740 14188 23792
rect 14240 23780 14246 23792
rect 15838 23780 15844 23792
rect 14240 23752 15844 23780
rect 14240 23740 14246 23752
rect 15838 23740 15844 23752
rect 15896 23740 15902 23792
rect 16853 23783 16911 23789
rect 16853 23749 16865 23783
rect 16899 23780 16911 23783
rect 17218 23780 17224 23792
rect 16899 23752 17224 23780
rect 16899 23749 16911 23752
rect 16853 23743 16911 23749
rect 17218 23740 17224 23752
rect 17276 23740 17282 23792
rect 18138 23740 18144 23792
rect 18196 23780 18202 23792
rect 18417 23783 18475 23789
rect 18417 23780 18429 23783
rect 18196 23752 18429 23780
rect 18196 23740 18202 23752
rect 18417 23749 18429 23752
rect 18463 23749 18475 23783
rect 18417 23743 18475 23749
rect 19886 23740 19892 23792
rect 19944 23740 19950 23792
rect 21358 23740 21364 23792
rect 21416 23780 21422 23792
rect 21818 23780 21824 23792
rect 21416 23752 21824 23780
rect 21416 23740 21422 23752
rect 21818 23740 21824 23752
rect 21876 23740 21882 23792
rect 25222 23740 25228 23792
rect 25280 23780 25286 23792
rect 29089 23783 29147 23789
rect 29089 23780 29101 23783
rect 25280 23752 29101 23780
rect 25280 23740 25286 23752
rect 29089 23749 29101 23752
rect 29135 23749 29147 23783
rect 29089 23743 29147 23749
rect 29270 23740 29276 23792
rect 29328 23740 29334 23792
rect 13357 23715 13415 23721
rect 13357 23681 13369 23715
rect 13403 23681 13415 23715
rect 13357 23675 13415 23681
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23681 13875 23715
rect 13817 23675 13875 23681
rect 12618 23604 12624 23656
rect 12676 23644 12682 23656
rect 13262 23644 13268 23656
rect 12676 23616 13268 23644
rect 12676 23604 12682 23616
rect 13262 23604 13268 23616
rect 13320 23604 13326 23656
rect 13832 23644 13860 23675
rect 13906 23672 13912 23724
rect 13964 23672 13970 23724
rect 14366 23721 14372 23724
rect 14323 23715 14372 23721
rect 14323 23681 14335 23715
rect 14369 23681 14372 23715
rect 14323 23675 14372 23681
rect 14366 23672 14372 23675
rect 14424 23672 14430 23724
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 14516 23684 15240 23712
rect 14516 23672 14522 23684
rect 15102 23644 15108 23656
rect 13832 23616 15108 23644
rect 15102 23604 15108 23616
rect 15160 23604 15166 23656
rect 15212 23644 15240 23684
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17494 23712 17500 23724
rect 17092 23684 17500 23712
rect 17092 23672 17098 23684
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 18877 23715 18935 23721
rect 18877 23712 18889 23715
rect 17604 23684 18889 23712
rect 17604 23644 17632 23684
rect 18877 23681 18889 23684
rect 18923 23681 18935 23715
rect 18877 23675 18935 23681
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19978 23672 19984 23724
rect 20036 23712 20042 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 20036 23684 20269 23712
rect 20036 23672 20042 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20257 23675 20315 23681
rect 20625 23715 20683 23721
rect 20625 23681 20637 23715
rect 20671 23712 20683 23715
rect 20898 23712 20904 23724
rect 20671 23684 20904 23712
rect 20671 23681 20683 23684
rect 20625 23675 20683 23681
rect 20898 23672 20904 23684
rect 20956 23712 20962 23724
rect 21174 23712 21180 23724
rect 20956 23684 21180 23712
rect 20956 23672 20962 23684
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 26786 23672 26792 23724
rect 26844 23672 26850 23724
rect 27154 23672 27160 23724
rect 27212 23672 27218 23724
rect 27430 23672 27436 23724
rect 27488 23672 27494 23724
rect 27522 23672 27528 23724
rect 27580 23712 27586 23724
rect 27801 23715 27859 23721
rect 27801 23712 27813 23715
rect 27580 23684 27813 23712
rect 27580 23672 27586 23684
rect 27801 23681 27813 23684
rect 27847 23681 27859 23715
rect 27801 23675 27859 23681
rect 28994 23672 29000 23724
rect 29052 23672 29058 23724
rect 15212 23616 17632 23644
rect 18785 23647 18843 23653
rect 18785 23613 18797 23647
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 10284 23548 12020 23576
rect 18800 23576 18828 23607
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 27249 23647 27307 23653
rect 19208 23616 21680 23644
rect 19208 23604 19214 23616
rect 20073 23579 20131 23585
rect 20073 23576 20085 23579
rect 18800 23548 20085 23576
rect 10284 23536 10290 23548
rect 20073 23545 20085 23548
rect 20119 23545 20131 23579
rect 20073 23539 20131 23545
rect 9766 23508 9772 23520
rect 7300 23480 9772 23508
rect 9766 23468 9772 23480
rect 9824 23508 9830 23520
rect 9950 23508 9956 23520
rect 9824 23480 9956 23508
rect 9824 23468 9830 23480
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10505 23511 10563 23517
rect 10505 23477 10517 23511
rect 10551 23508 10563 23511
rect 11054 23508 11060 23520
rect 10551 23480 11060 23508
rect 10551 23477 10563 23480
rect 10505 23471 10563 23477
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 11149 23511 11207 23517
rect 11149 23477 11161 23511
rect 11195 23508 11207 23511
rect 11238 23508 11244 23520
rect 11195 23480 11244 23508
rect 11195 23477 11207 23480
rect 11149 23471 11207 23477
rect 11238 23468 11244 23480
rect 11296 23468 11302 23520
rect 13449 23511 13507 23517
rect 13449 23477 13461 23511
rect 13495 23508 13507 23511
rect 13538 23508 13544 23520
rect 13495 23480 13544 23508
rect 13495 23477 13507 23480
rect 13449 23471 13507 23477
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 16669 23511 16727 23517
rect 16669 23477 16681 23511
rect 16715 23508 16727 23511
rect 16850 23508 16856 23520
rect 16715 23480 16856 23508
rect 16715 23477 16727 23480
rect 16669 23471 16727 23477
rect 16850 23468 16856 23480
rect 16908 23468 16914 23520
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 17000 23480 18521 23508
rect 17000 23468 17006 23480
rect 18509 23477 18521 23480
rect 18555 23508 18567 23511
rect 18874 23508 18880 23520
rect 18555 23480 18880 23508
rect 18555 23477 18567 23480
rect 18509 23471 18567 23477
rect 18874 23468 18880 23480
rect 18932 23468 18938 23520
rect 19061 23511 19119 23517
rect 19061 23477 19073 23511
rect 19107 23508 19119 23511
rect 19794 23508 19800 23520
rect 19107 23480 19800 23508
rect 19107 23477 19119 23480
rect 19061 23471 19119 23477
rect 19794 23468 19800 23480
rect 19852 23468 19858 23520
rect 19886 23468 19892 23520
rect 19944 23468 19950 23520
rect 20530 23468 20536 23520
rect 20588 23508 20594 23520
rect 21542 23508 21548 23520
rect 20588 23480 21548 23508
rect 20588 23468 20594 23480
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 21652 23508 21680 23616
rect 27249 23613 27261 23647
rect 27295 23613 27307 23647
rect 27249 23607 27307 23613
rect 26513 23579 26571 23585
rect 26513 23545 26525 23579
rect 26559 23576 26571 23579
rect 26973 23579 27031 23585
rect 26973 23576 26985 23579
rect 26559 23548 26985 23576
rect 26559 23545 26571 23548
rect 26513 23539 26571 23545
rect 26973 23545 26985 23548
rect 27019 23545 27031 23579
rect 27264 23576 27292 23607
rect 27338 23604 27344 23656
rect 27396 23604 27402 23656
rect 27540 23576 27568 23672
rect 27706 23604 27712 23656
rect 27764 23604 27770 23656
rect 27264 23548 27568 23576
rect 26973 23539 27031 23545
rect 27890 23508 27896 23520
rect 21652 23480 27896 23508
rect 27890 23468 27896 23480
rect 27948 23468 27954 23520
rect 1104 23418 29716 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 29716 23418
rect 1104 23344 29716 23366
rect 4433 23307 4491 23313
rect 4433 23273 4445 23307
rect 4479 23304 4491 23307
rect 4614 23304 4620 23316
rect 4479 23276 4620 23304
rect 4479 23273 4491 23276
rect 4433 23267 4491 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 5905 23307 5963 23313
rect 5905 23304 5917 23307
rect 5684 23276 5917 23304
rect 5684 23264 5690 23276
rect 5905 23273 5917 23276
rect 5951 23273 5963 23307
rect 5905 23267 5963 23273
rect 8021 23307 8079 23313
rect 8021 23273 8033 23307
rect 8067 23304 8079 23307
rect 11238 23304 11244 23316
rect 8067 23276 11244 23304
rect 8067 23273 8079 23276
rect 8021 23267 8079 23273
rect 11238 23264 11244 23276
rect 11296 23264 11302 23316
rect 12250 23264 12256 23316
rect 12308 23264 12314 23316
rect 12897 23307 12955 23313
rect 12897 23273 12909 23307
rect 12943 23304 12955 23307
rect 12986 23304 12992 23316
rect 12943 23276 12992 23304
rect 12943 23273 12955 23276
rect 12897 23267 12955 23273
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 15565 23307 15623 23313
rect 14936 23276 15148 23304
rect 7190 23196 7196 23248
rect 7248 23236 7254 23248
rect 8205 23239 8263 23245
rect 8205 23236 8217 23239
rect 7248 23208 8217 23236
rect 7248 23196 7254 23208
rect 8205 23205 8217 23208
rect 8251 23205 8263 23239
rect 8205 23199 8263 23205
rect 9766 23196 9772 23248
rect 9824 23236 9830 23248
rect 10594 23236 10600 23248
rect 9824 23208 10600 23236
rect 9824 23196 9830 23208
rect 10594 23196 10600 23208
rect 10652 23236 10658 23248
rect 12713 23239 12771 23245
rect 10652 23208 12572 23236
rect 10652 23196 10658 23208
rect 4430 23168 4436 23180
rect 4356 23140 4436 23168
rect 4356 23109 4384 23140
rect 4430 23128 4436 23140
rect 4488 23168 4494 23180
rect 4488 23140 5396 23168
rect 4488 23128 4494 23140
rect 5368 23112 5396 23140
rect 9306 23128 9312 23180
rect 9364 23168 9370 23180
rect 10870 23168 10876 23180
rect 9364 23140 10876 23168
rect 9364 23128 9370 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 12434 23128 12440 23180
rect 12492 23128 12498 23180
rect 12544 23168 12572 23208
rect 12713 23205 12725 23239
rect 12759 23236 12771 23239
rect 13906 23236 13912 23248
rect 12759 23208 13912 23236
rect 12759 23205 12771 23208
rect 12713 23199 12771 23205
rect 13906 23196 13912 23208
rect 13964 23196 13970 23248
rect 14090 23196 14096 23248
rect 14148 23236 14154 23248
rect 14148 23208 14504 23236
rect 14148 23196 14154 23208
rect 12544 23140 12848 23168
rect 4341 23103 4399 23109
rect 4341 23069 4353 23103
rect 4387 23069 4399 23103
rect 4341 23063 4399 23069
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23100 4583 23103
rect 4798 23100 4804 23112
rect 4571 23072 4804 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 4798 23060 4804 23072
rect 4856 23060 4862 23112
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 5718 23060 5724 23112
rect 5776 23060 5782 23112
rect 7374 23060 7380 23112
rect 7432 23060 7438 23112
rect 7466 23060 7472 23112
rect 7524 23100 7530 23112
rect 7883 23103 7941 23109
rect 7524 23072 7569 23100
rect 7524 23060 7530 23072
rect 7883 23069 7895 23103
rect 7929 23100 7941 23103
rect 8018 23100 8024 23112
rect 7929 23072 8024 23100
rect 7929 23069 7941 23072
rect 7883 23063 7941 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 8297 23103 8355 23109
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 10042 23100 10048 23112
rect 8343 23072 10048 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 10226 23060 10232 23112
rect 10284 23100 10290 23112
rect 10965 23103 11023 23109
rect 10965 23100 10977 23103
rect 10284 23072 10977 23100
rect 10284 23060 10290 23072
rect 10965 23069 10977 23072
rect 11011 23069 11023 23103
rect 10965 23063 11023 23069
rect 11054 23060 11060 23112
rect 11112 23060 11118 23112
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 12820 23109 12848 23140
rect 14366 23128 14372 23180
rect 14424 23128 14430 23180
rect 12529 23103 12587 23109
rect 11296 23072 12434 23100
rect 11296 23060 11302 23072
rect 2682 22992 2688 23044
rect 2740 23032 2746 23044
rect 5258 23032 5264 23044
rect 2740 23004 5264 23032
rect 2740 22992 2746 23004
rect 5258 22992 5264 23004
rect 5316 22992 5322 23044
rect 5534 22992 5540 23044
rect 5592 22992 5598 23044
rect 5629 23035 5687 23041
rect 5629 23001 5641 23035
rect 5675 23001 5687 23035
rect 5629 22995 5687 23001
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 5644 22964 5672 22995
rect 7650 22992 7656 23044
rect 7708 22992 7714 23044
rect 7745 23035 7803 23041
rect 7745 23001 7757 23035
rect 7791 23001 7803 23035
rect 7745 22995 7803 23001
rect 11333 23035 11391 23041
rect 11333 23001 11345 23035
rect 11379 23032 11391 23035
rect 12253 23035 12311 23041
rect 12253 23032 12265 23035
rect 11379 23004 12265 23032
rect 11379 23001 11391 23004
rect 11333 22995 11391 23001
rect 12253 23001 12265 23004
rect 12299 23001 12311 23035
rect 12406 23032 12434 23072
rect 12529 23069 12541 23103
rect 12575 23069 12587 23103
rect 12529 23063 12587 23069
rect 12805 23103 12863 23109
rect 12805 23069 12817 23103
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 12544 23032 12572 23063
rect 14090 23060 14096 23112
rect 14148 23060 14154 23112
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23100 14243 23103
rect 14274 23100 14280 23112
rect 14231 23072 14280 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 14476 23109 14504 23208
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14829 23103 14887 23109
rect 14829 23069 14841 23103
rect 14875 23100 14887 23103
rect 14936 23100 14964 23276
rect 15013 23239 15071 23245
rect 15013 23205 15025 23239
rect 15059 23205 15071 23239
rect 15120 23236 15148 23276
rect 15565 23273 15577 23307
rect 15611 23304 15623 23307
rect 16117 23307 16175 23313
rect 16117 23304 16129 23307
rect 15611 23276 16129 23304
rect 15611 23273 15623 23276
rect 15565 23267 15623 23273
rect 16117 23273 16129 23276
rect 16163 23273 16175 23307
rect 16117 23267 16175 23273
rect 16577 23307 16635 23313
rect 16577 23273 16589 23307
rect 16623 23304 16635 23307
rect 16666 23304 16672 23316
rect 16623 23276 16672 23304
rect 16623 23273 16635 23276
rect 16577 23267 16635 23273
rect 16666 23264 16672 23276
rect 16724 23304 16730 23316
rect 16942 23304 16948 23316
rect 16724 23276 16948 23304
rect 16724 23264 16730 23276
rect 16942 23264 16948 23276
rect 17000 23264 17006 23316
rect 18322 23264 18328 23316
rect 18380 23304 18386 23316
rect 18969 23307 19027 23313
rect 18969 23304 18981 23307
rect 18380 23276 18981 23304
rect 18380 23264 18386 23276
rect 18969 23273 18981 23276
rect 19015 23304 19027 23307
rect 19150 23304 19156 23316
rect 19015 23276 19156 23304
rect 19015 23273 19027 23276
rect 18969 23267 19027 23273
rect 19150 23264 19156 23276
rect 19208 23264 19214 23316
rect 21726 23264 21732 23316
rect 21784 23264 21790 23316
rect 27249 23307 27307 23313
rect 27249 23273 27261 23307
rect 27295 23304 27307 23307
rect 27706 23304 27712 23316
rect 27295 23276 27712 23304
rect 27295 23273 27307 23276
rect 27249 23267 27307 23273
rect 27706 23264 27712 23276
rect 27764 23304 27770 23316
rect 27764 23276 28304 23304
rect 27764 23264 27770 23276
rect 15194 23236 15200 23248
rect 15120 23208 15200 23236
rect 15013 23199 15071 23205
rect 14875 23072 14964 23100
rect 15028 23100 15056 23199
rect 15194 23196 15200 23208
rect 15252 23236 15258 23248
rect 15841 23239 15899 23245
rect 15841 23236 15853 23239
rect 15252 23208 15853 23236
rect 15252 23196 15258 23208
rect 15841 23205 15853 23208
rect 15887 23205 15899 23239
rect 17037 23239 17095 23245
rect 15841 23199 15899 23205
rect 16408 23208 16896 23236
rect 15657 23171 15715 23177
rect 15657 23168 15669 23171
rect 15304 23140 15669 23168
rect 15304 23109 15332 23140
rect 15657 23137 15669 23140
rect 15703 23137 15715 23171
rect 15657 23131 15715 23137
rect 16408 23112 16436 23208
rect 15289 23103 15347 23109
rect 15289 23100 15301 23103
rect 15028 23072 15301 23100
rect 14875 23069 14887 23072
rect 14829 23063 14887 23069
rect 15289 23069 15301 23072
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 15378 23060 15384 23112
rect 15436 23060 15442 23112
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 15933 23103 15991 23109
rect 15933 23100 15945 23103
rect 15528 23072 15945 23100
rect 15528 23060 15534 23072
rect 15933 23069 15945 23072
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 16390 23060 16396 23112
rect 16448 23060 16454 23112
rect 16666 23060 16672 23112
rect 16724 23060 16730 23112
rect 16761 23103 16819 23109
rect 16761 23069 16773 23103
rect 16807 23069 16819 23103
rect 16868 23100 16896 23208
rect 17037 23205 17049 23239
rect 17083 23205 17095 23239
rect 17037 23199 17095 23205
rect 17313 23239 17371 23245
rect 17313 23205 17325 23239
rect 17359 23236 17371 23239
rect 17359 23208 18828 23236
rect 17359 23205 17371 23208
rect 17313 23199 17371 23205
rect 17052 23168 17080 23199
rect 17052 23140 17356 23168
rect 17328 23109 17356 23140
rect 17697 23140 18184 23168
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16868 23072 17141 23100
rect 16761 23063 16819 23069
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 17313 23103 17371 23109
rect 17313 23069 17325 23103
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 12406 23004 12572 23032
rect 14292 23032 14320 23060
rect 14645 23035 14703 23041
rect 14645 23032 14657 23035
rect 14292 23004 14657 23032
rect 12253 22995 12311 23001
rect 14645 23001 14657 23004
rect 14691 23001 14703 23035
rect 14645 22995 14703 23001
rect 7760 22964 7788 22995
rect 14734 22992 14740 23044
rect 14792 22992 14798 23044
rect 15565 23035 15623 23041
rect 15565 23032 15577 23035
rect 14936 23004 15577 23032
rect 4948 22936 7788 22964
rect 14369 22967 14427 22973
rect 4948 22924 4954 22936
rect 14369 22933 14381 22967
rect 14415 22964 14427 22967
rect 14936 22964 14964 23004
rect 15565 23001 15577 23004
rect 15611 23001 15623 23035
rect 15565 22995 15623 23001
rect 15657 23035 15715 23041
rect 15657 23001 15669 23035
rect 15703 23032 15715 23035
rect 16776 23032 16804 23063
rect 15703 23004 16804 23032
rect 15703 23001 15715 23004
rect 15657 22995 15715 23001
rect 16850 22992 16856 23044
rect 16908 22992 16914 23044
rect 16942 22992 16948 23044
rect 17000 23032 17006 23044
rect 17037 23035 17095 23041
rect 17037 23032 17049 23035
rect 17000 23004 17049 23032
rect 17000 22992 17006 23004
rect 17037 23001 17049 23004
rect 17083 23001 17095 23035
rect 17037 22995 17095 23001
rect 14415 22936 14964 22964
rect 14415 22933 14427 22936
rect 14369 22927 14427 22933
rect 15102 22924 15108 22976
rect 15160 22924 15166 22976
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 17697 22964 17725 23140
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23069 17831 23103
rect 17773 23063 17831 23069
rect 17788 23032 17816 23063
rect 17954 23060 17960 23112
rect 18012 23060 18018 23112
rect 18046 23060 18052 23112
rect 18104 23060 18110 23112
rect 18156 23109 18184 23140
rect 18141 23103 18199 23109
rect 18141 23069 18153 23103
rect 18187 23100 18199 23103
rect 18322 23100 18328 23112
rect 18187 23072 18328 23100
rect 18187 23069 18199 23072
rect 18141 23063 18199 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 18690 23060 18696 23112
rect 18748 23060 18754 23112
rect 18800 23109 18828 23208
rect 19058 23196 19064 23248
rect 19116 23236 19122 23248
rect 19116 23208 22094 23236
rect 19116 23196 19122 23208
rect 22066 23168 22094 23208
rect 23842 23196 23848 23248
rect 23900 23236 23906 23248
rect 23900 23208 24808 23236
rect 23900 23196 23906 23208
rect 23566 23168 23572 23180
rect 22066 23140 23572 23168
rect 23566 23128 23572 23140
rect 23624 23168 23630 23180
rect 24673 23171 24731 23177
rect 24673 23168 24685 23171
rect 23624 23140 24685 23168
rect 23624 23128 23630 23140
rect 24673 23137 24685 23140
rect 24719 23137 24731 23171
rect 24673 23131 24731 23137
rect 18785 23103 18843 23109
rect 18785 23069 18797 23103
rect 18831 23069 18843 23103
rect 18785 23063 18843 23069
rect 19061 23103 19119 23109
rect 19061 23069 19073 23103
rect 19107 23100 19119 23103
rect 19426 23100 19432 23112
rect 19107 23072 19432 23100
rect 19107 23069 19119 23072
rect 19061 23063 19119 23069
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23100 21327 23103
rect 21726 23100 21732 23112
rect 21315 23072 21732 23100
rect 21315 23069 21327 23072
rect 21269 23063 21327 23069
rect 21726 23060 21732 23072
rect 21784 23060 21790 23112
rect 24489 23103 24547 23109
rect 24489 23069 24501 23103
rect 24535 23069 24547 23103
rect 24489 23063 24547 23069
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24780 23100 24808 23208
rect 24857 23171 24915 23177
rect 24857 23137 24869 23171
rect 24903 23168 24915 23171
rect 28166 23168 28172 23180
rect 24903 23140 28172 23168
rect 24903 23137 24915 23140
rect 24857 23131 24915 23137
rect 28166 23128 28172 23140
rect 28224 23128 28230 23180
rect 28276 23177 28304 23276
rect 28261 23171 28319 23177
rect 28261 23137 28273 23171
rect 28307 23137 28319 23171
rect 28261 23131 28319 23137
rect 24627 23072 24808 23100
rect 25133 23103 25191 23109
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 25133 23069 25145 23103
rect 25179 23100 25191 23103
rect 26234 23100 26240 23112
rect 25179 23072 26240 23100
rect 25179 23069 25191 23072
rect 25133 23063 25191 23069
rect 18509 23035 18567 23041
rect 18509 23032 18521 23035
rect 17788 23004 18521 23032
rect 18509 23001 18521 23004
rect 18555 23001 18567 23035
rect 18509 22995 18567 23001
rect 23201 23035 23259 23041
rect 23201 23001 23213 23035
rect 23247 23032 23259 23035
rect 23658 23032 23664 23044
rect 23247 23004 23664 23032
rect 23247 23001 23259 23004
rect 23201 22995 23259 23001
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 24504 23032 24532 23063
rect 26234 23060 26240 23072
rect 26292 23060 26298 23112
rect 27154 23060 27160 23112
rect 27212 23060 27218 23112
rect 27338 23060 27344 23112
rect 27396 23100 27402 23112
rect 27801 23103 27859 23109
rect 27396 23072 27660 23100
rect 27396 23060 27402 23072
rect 25406 23032 25412 23044
rect 24504 23004 25412 23032
rect 25406 22992 25412 23004
rect 25464 22992 25470 23044
rect 27172 23032 27200 23060
rect 27632 23041 27660 23072
rect 27801 23069 27813 23103
rect 27847 23100 27859 23103
rect 28077 23103 28135 23109
rect 28077 23100 28089 23103
rect 27847 23072 28089 23100
rect 27847 23069 27859 23072
rect 27801 23063 27859 23069
rect 28077 23069 28089 23072
rect 28123 23069 28135 23103
rect 28077 23063 28135 23069
rect 27433 23035 27491 23041
rect 27433 23032 27445 23035
rect 27172 23004 27445 23032
rect 27433 23001 27445 23004
rect 27479 23001 27491 23035
rect 27433 22995 27491 23001
rect 27617 23035 27675 23041
rect 27617 23001 27629 23035
rect 27663 23032 27675 23035
rect 27706 23032 27712 23044
rect 27663 23004 27712 23032
rect 27663 23001 27675 23004
rect 27617 22995 27675 23001
rect 27706 22992 27712 23004
rect 27764 22992 27770 23044
rect 16724 22936 17725 22964
rect 18417 22967 18475 22973
rect 16724 22924 16730 22936
rect 18417 22933 18429 22967
rect 18463 22964 18475 22967
rect 20438 22964 20444 22976
rect 18463 22936 20444 22964
rect 18463 22933 18475 22936
rect 18417 22927 18475 22933
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 21450 22924 21456 22976
rect 21508 22964 21514 22976
rect 21818 22964 21824 22976
rect 21508 22936 21824 22964
rect 21508 22924 21514 22936
rect 21818 22924 21824 22936
rect 21876 22964 21882 22976
rect 22002 22964 22008 22976
rect 21876 22936 22008 22964
rect 21876 22924 21882 22936
rect 22002 22924 22008 22936
rect 22060 22924 22066 22976
rect 25038 22924 25044 22976
rect 25096 22924 25102 22976
rect 27890 22924 27896 22976
rect 27948 22924 27954 22976
rect 1104 22874 29716 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 29716 22874
rect 1104 22800 29716 22822
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 4525 22763 4583 22769
rect 4525 22760 4537 22763
rect 4488 22732 4537 22760
rect 4488 22720 4494 22732
rect 4525 22729 4537 22732
rect 4571 22729 4583 22763
rect 4525 22723 4583 22729
rect 5368 22732 7926 22760
rect 1673 22627 1731 22633
rect 1673 22593 1685 22627
rect 1719 22624 1731 22627
rect 2682 22624 2688 22636
rect 1719 22596 2688 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 2682 22584 2688 22596
rect 2740 22584 2746 22636
rect 2774 22584 2780 22636
rect 2832 22584 2838 22636
rect 4154 22584 4160 22636
rect 4212 22584 4218 22636
rect 4540 22624 4568 22723
rect 4798 22652 4804 22704
rect 4856 22692 4862 22704
rect 5077 22695 5135 22701
rect 5077 22692 5089 22695
rect 4856 22664 5089 22692
rect 4856 22652 4862 22664
rect 5077 22661 5089 22664
rect 5123 22661 5135 22695
rect 5077 22655 5135 22661
rect 5368 22633 5396 22732
rect 5534 22652 5540 22704
rect 5592 22692 5598 22704
rect 6089 22695 6147 22701
rect 6089 22692 6101 22695
rect 5592 22664 6101 22692
rect 5592 22652 5598 22664
rect 6089 22661 6101 22664
rect 6135 22661 6147 22695
rect 6730 22692 6736 22704
rect 6089 22655 6147 22661
rect 6288 22664 6736 22692
rect 4893 22627 4951 22633
rect 4893 22624 4905 22627
rect 4540 22596 4905 22624
rect 4893 22593 4905 22596
rect 4939 22593 4951 22627
rect 4893 22587 4951 22593
rect 5353 22627 5411 22633
rect 5353 22593 5365 22627
rect 5399 22593 5411 22627
rect 5353 22587 5411 22593
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22593 5687 22627
rect 5629 22587 5687 22593
rect 842 22516 848 22568
rect 900 22556 906 22568
rect 1397 22559 1455 22565
rect 1397 22556 1409 22559
rect 900 22528 1409 22556
rect 900 22516 906 22528
rect 1397 22525 1409 22528
rect 1443 22525 1455 22559
rect 1397 22519 1455 22525
rect 3050 22516 3056 22568
rect 3108 22516 3114 22568
rect 5644 22488 5672 22587
rect 5718 22584 5724 22636
rect 5776 22584 5782 22636
rect 6181 22627 6239 22633
rect 6181 22593 6193 22627
rect 6227 22624 6239 22627
rect 6288 22624 6316 22664
rect 6730 22652 6736 22664
rect 6788 22652 6794 22704
rect 6914 22652 6920 22704
rect 6972 22692 6978 22704
rect 7650 22692 7656 22704
rect 6972 22664 7656 22692
rect 6972 22652 6978 22664
rect 7650 22652 7656 22664
rect 7708 22652 7714 22704
rect 6227 22596 6316 22624
rect 6227 22593 6239 22596
rect 6181 22587 6239 22593
rect 6362 22584 6368 22636
rect 6420 22584 6426 22636
rect 7537 22627 7595 22633
rect 7537 22593 7549 22627
rect 7583 22624 7595 22627
rect 7583 22622 7604 22624
rect 7583 22594 7696 22622
rect 7583 22593 7595 22594
rect 7537 22587 7595 22593
rect 5736 22556 5764 22584
rect 6457 22559 6515 22565
rect 6457 22556 6469 22559
rect 5736 22528 6469 22556
rect 6457 22525 6469 22528
rect 6503 22525 6515 22559
rect 6457 22519 6515 22525
rect 6546 22516 6552 22568
rect 6604 22556 6610 22568
rect 7668 22556 7696 22594
rect 7742 22584 7748 22636
rect 7800 22584 7806 22636
rect 7898 22633 7926 22732
rect 8018 22720 8024 22772
rect 8076 22760 8082 22772
rect 8202 22760 8208 22772
rect 8076 22732 8208 22760
rect 8076 22720 8082 22732
rect 8202 22720 8208 22732
rect 8260 22760 8266 22772
rect 9033 22763 9091 22769
rect 9033 22760 9045 22763
rect 8260 22732 9045 22760
rect 8260 22720 8266 22732
rect 9033 22729 9045 22732
rect 9079 22729 9091 22763
rect 9033 22723 9091 22729
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 9732 22732 9873 22760
rect 9732 22720 9738 22732
rect 9861 22729 9873 22732
rect 9907 22760 9919 22763
rect 9950 22760 9956 22772
rect 9907 22732 9956 22760
rect 9907 22729 9919 22732
rect 9861 22723 9919 22729
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 10870 22720 10876 22772
rect 10928 22720 10934 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15470 22760 15476 22772
rect 14792 22732 15476 22760
rect 14792 22720 14798 22732
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 16448 22732 16681 22760
rect 16448 22720 16454 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 17402 22760 17408 22772
rect 16669 22723 16727 22729
rect 17236 22732 17408 22760
rect 10505 22695 10563 22701
rect 10505 22692 10517 22695
rect 8312 22664 10517 22692
rect 7883 22627 7941 22633
rect 7883 22593 7895 22627
rect 7929 22624 7941 22627
rect 8110 22624 8116 22636
rect 7929 22596 8116 22624
rect 7929 22593 7941 22596
rect 7883 22587 7941 22593
rect 8110 22584 8116 22596
rect 8168 22584 8174 22636
rect 8202 22556 8208 22568
rect 6604 22528 7512 22556
rect 7668 22528 8208 22556
rect 6604 22516 6610 22528
rect 6178 22488 6184 22500
rect 5644 22460 6184 22488
rect 6178 22448 6184 22460
rect 6236 22488 6242 22500
rect 6914 22488 6920 22500
rect 6236 22460 6920 22488
rect 6236 22448 6242 22460
rect 6914 22448 6920 22460
rect 6972 22448 6978 22500
rect 4706 22380 4712 22432
rect 4764 22380 4770 22432
rect 5626 22380 5632 22432
rect 5684 22420 5690 22432
rect 5905 22423 5963 22429
rect 5905 22420 5917 22423
rect 5684 22392 5917 22420
rect 5684 22380 5690 22392
rect 5905 22389 5917 22392
rect 5951 22389 5963 22423
rect 5905 22383 5963 22389
rect 7374 22380 7380 22432
rect 7432 22380 7438 22432
rect 7484 22420 7512 22528
rect 8202 22516 8208 22528
rect 8260 22516 8266 22568
rect 7742 22448 7748 22500
rect 7800 22488 7806 22500
rect 8312 22488 8340 22664
rect 10505 22661 10517 22664
rect 10551 22661 10563 22695
rect 10888 22692 10916 22720
rect 10888 22664 11008 22692
rect 10505 22655 10563 22661
rect 8938 22584 8944 22636
rect 8996 22624 9002 22636
rect 9125 22627 9183 22633
rect 9125 22624 9137 22627
rect 8996 22596 9137 22624
rect 8996 22584 9002 22596
rect 9125 22593 9137 22596
rect 9171 22593 9183 22627
rect 9125 22587 9183 22593
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22624 10011 22627
rect 10318 22624 10324 22636
rect 9999 22596 10324 22624
rect 9999 22593 10011 22596
rect 9953 22587 10011 22593
rect 9140 22556 9168 22587
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 10781 22627 10839 22633
rect 10781 22593 10793 22627
rect 10827 22624 10839 22627
rect 10870 22624 10876 22636
rect 10827 22596 10876 22624
rect 10827 22593 10839 22596
rect 10781 22587 10839 22593
rect 10502 22556 10508 22568
rect 9140 22528 10508 22556
rect 10502 22516 10508 22528
rect 10560 22516 10566 22568
rect 10612 22556 10640 22587
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 10980 22633 11008 22664
rect 12986 22652 12992 22704
rect 13044 22652 13050 22704
rect 14366 22652 14372 22704
rect 14424 22692 14430 22704
rect 16850 22692 16856 22704
rect 14424 22664 16856 22692
rect 14424 22652 14430 22664
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 17236 22701 17264 22732
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 18046 22760 18052 22772
rect 17696 22732 18052 22760
rect 17221 22695 17279 22701
rect 17221 22661 17233 22695
rect 17267 22661 17279 22695
rect 17221 22655 17279 22661
rect 17310 22652 17316 22704
rect 17368 22652 17374 22704
rect 17696 22692 17724 22732
rect 18046 22720 18052 22732
rect 18104 22760 18110 22772
rect 18969 22763 19027 22769
rect 18969 22760 18981 22763
rect 18104 22732 18981 22760
rect 18104 22720 18110 22732
rect 18969 22729 18981 22732
rect 19015 22729 19027 22763
rect 19702 22760 19708 22772
rect 18969 22723 19027 22729
rect 19076 22732 19708 22760
rect 17604 22664 17724 22692
rect 17865 22695 17923 22701
rect 10965 22627 11023 22633
rect 10965 22593 10977 22627
rect 11011 22624 11023 22627
rect 11609 22627 11667 22633
rect 11609 22624 11621 22627
rect 11011 22596 11621 22624
rect 11011 22593 11023 22596
rect 10965 22587 11023 22593
rect 11609 22593 11621 22596
rect 11655 22593 11667 22627
rect 11609 22587 11667 22593
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22593 12863 22627
rect 12805 22587 12863 22593
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22624 13231 22627
rect 13262 22624 13268 22636
rect 13219 22596 13268 22624
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 12158 22556 12164 22568
rect 10612 22528 12164 22556
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12710 22556 12716 22568
rect 12406 22528 12716 22556
rect 12406 22488 12434 22528
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 7800 22460 8340 22488
rect 10704 22460 12434 22488
rect 12820 22488 12848 22587
rect 12912 22556 12940 22587
rect 13262 22584 13268 22596
rect 13320 22584 13326 22636
rect 16114 22584 16120 22636
rect 16172 22624 16178 22636
rect 16942 22624 16948 22636
rect 16172 22596 16948 22624
rect 16172 22584 16178 22596
rect 16942 22584 16948 22596
rect 17000 22584 17006 22636
rect 17604 22633 17632 22664
rect 17865 22661 17877 22695
rect 17911 22661 17923 22695
rect 17865 22655 17923 22661
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22593 17647 22627
rect 17589 22587 17647 22593
rect 17678 22584 17684 22636
rect 17736 22584 17742 22636
rect 13722 22556 13728 22568
rect 12912 22528 13728 22556
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 16853 22559 16911 22565
rect 16853 22525 16865 22559
rect 16899 22556 16911 22559
rect 17697 22556 17725 22584
rect 17880 22568 17908 22655
rect 17954 22652 17960 22704
rect 18012 22652 18018 22704
rect 18322 22652 18328 22704
rect 18380 22652 18386 22704
rect 16899 22528 17725 22556
rect 16899 22525 16911 22528
rect 16853 22519 16911 22525
rect 17862 22516 17868 22568
rect 17920 22516 17926 22568
rect 17972 22556 18000 22652
rect 18095 22627 18153 22633
rect 18095 22593 18107 22627
rect 18141 22624 18153 22627
rect 18414 22624 18420 22636
rect 18141 22596 18420 22624
rect 18141 22593 18153 22596
rect 18095 22587 18153 22593
rect 18414 22584 18420 22596
rect 18472 22624 18478 22636
rect 18509 22627 18567 22633
rect 18509 22624 18521 22627
rect 18472 22596 18521 22624
rect 18472 22584 18478 22596
rect 18509 22593 18521 22596
rect 18555 22593 18567 22627
rect 18509 22587 18567 22593
rect 18601 22627 18659 22633
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18877 22627 18935 22633
rect 18877 22593 18889 22627
rect 18923 22624 18935 22627
rect 19076 22624 19104 22732
rect 19702 22720 19708 22732
rect 19760 22760 19766 22772
rect 19760 22732 20668 22760
rect 19760 22720 19766 22732
rect 19245 22695 19303 22701
rect 19245 22661 19257 22695
rect 19291 22692 19303 22695
rect 19426 22692 19432 22704
rect 19291 22664 19432 22692
rect 19291 22661 19303 22664
rect 19245 22655 19303 22661
rect 19426 22652 19432 22664
rect 19484 22692 19490 22704
rect 20162 22692 20168 22704
rect 19484 22664 20168 22692
rect 19484 22652 19490 22664
rect 20162 22652 20168 22664
rect 20220 22692 20226 22704
rect 20220 22664 20392 22692
rect 20220 22652 20226 22664
rect 18923 22596 19104 22624
rect 18923 22593 18935 22596
rect 18877 22587 18935 22593
rect 18616 22556 18644 22587
rect 19150 22584 19156 22636
rect 19208 22584 19214 22636
rect 19337 22627 19395 22633
rect 19337 22593 19349 22627
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22624 19579 22627
rect 19702 22624 19708 22636
rect 19567 22596 19708 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 17972 22528 18644 22556
rect 18785 22559 18843 22565
rect 18785 22525 18797 22559
rect 18831 22556 18843 22559
rect 19352 22556 19380 22587
rect 19702 22584 19708 22596
rect 19760 22584 19766 22636
rect 19794 22584 19800 22636
rect 19852 22584 19858 22636
rect 19978 22584 19984 22636
rect 20036 22584 20042 22636
rect 20364 22633 20392 22664
rect 20640 22633 20668 22732
rect 21174 22720 21180 22772
rect 21232 22720 21238 22772
rect 21726 22720 21732 22772
rect 21784 22760 21790 22772
rect 23382 22760 23388 22772
rect 21784 22732 23388 22760
rect 21784 22720 21790 22732
rect 23382 22720 23388 22732
rect 23440 22760 23446 22772
rect 23440 22732 23704 22760
rect 23440 22720 23446 22732
rect 21545 22695 21603 22701
rect 21545 22661 21557 22695
rect 21591 22692 21603 22695
rect 21591 22664 22586 22692
rect 21591 22661 21603 22664
rect 21545 22655 21603 22661
rect 20349 22627 20407 22633
rect 20349 22593 20361 22627
rect 20395 22593 20407 22627
rect 20349 22587 20407 22593
rect 20625 22627 20683 22633
rect 20625 22593 20637 22627
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 20714 22584 20720 22636
rect 20772 22624 20778 22636
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20772 22596 20913 22624
rect 20772 22584 20778 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 20990 22584 20996 22636
rect 21048 22584 21054 22636
rect 21450 22584 21456 22636
rect 21508 22584 21514 22636
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 23676 22633 23704 22732
rect 25406 22720 25412 22772
rect 25464 22720 25470 22772
rect 27706 22720 27712 22772
rect 27764 22760 27770 22772
rect 29365 22763 29423 22769
rect 29365 22760 29377 22763
rect 27764 22732 29377 22760
rect 27764 22720 27770 22732
rect 29365 22729 29377 22732
rect 29411 22729 29423 22763
rect 29365 22723 29423 22729
rect 23934 22652 23940 22704
rect 23992 22652 23998 22704
rect 27890 22652 27896 22704
rect 27948 22652 27954 22704
rect 28902 22652 28908 22704
rect 28960 22652 28966 22704
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21784 22596 21833 22624
rect 21784 22584 21790 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 23661 22627 23719 22633
rect 23661 22593 23673 22627
rect 23707 22593 23719 22627
rect 23661 22587 23719 22593
rect 25038 22584 25044 22636
rect 25096 22584 25102 22636
rect 26234 22584 26240 22636
rect 26292 22624 26298 22636
rect 27157 22627 27215 22633
rect 27157 22624 27169 22627
rect 26292 22596 27169 22624
rect 26292 22584 26298 22596
rect 27157 22593 27169 22596
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 18831 22528 19380 22556
rect 18831 22525 18843 22528
rect 18785 22519 18843 22525
rect 18892 22500 18920 22528
rect 19886 22516 19892 22568
rect 19944 22556 19950 22568
rect 20073 22559 20131 22565
rect 20073 22556 20085 22559
rect 19944 22528 20085 22556
rect 19944 22516 19950 22528
rect 20073 22525 20085 22528
rect 20119 22525 20131 22559
rect 20073 22519 20131 22525
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22556 20223 22559
rect 20254 22556 20260 22568
rect 20211 22528 20260 22556
rect 20211 22525 20223 22528
rect 20165 22519 20223 22525
rect 20254 22516 20260 22528
rect 20312 22516 20318 22568
rect 20438 22516 20444 22568
rect 20496 22556 20502 22568
rect 22097 22559 22155 22565
rect 22097 22556 22109 22559
rect 20496 22528 22109 22556
rect 20496 22516 20502 22528
rect 22097 22525 22109 22528
rect 22143 22525 22155 22559
rect 22097 22519 22155 22525
rect 27614 22516 27620 22568
rect 27672 22516 27678 22568
rect 13538 22488 13544 22500
rect 12820 22460 13544 22488
rect 7800 22448 7806 22460
rect 10704 22420 10732 22460
rect 13538 22448 13544 22460
rect 13596 22448 13602 22500
rect 14734 22448 14740 22500
rect 14792 22488 14798 22500
rect 14918 22488 14924 22500
rect 14792 22460 14924 22488
rect 14792 22448 14798 22460
rect 14918 22448 14924 22460
rect 14976 22448 14982 22500
rect 15378 22448 15384 22500
rect 15436 22488 15442 22500
rect 18233 22491 18291 22497
rect 18233 22488 18245 22491
rect 15436 22460 18245 22488
rect 15436 22448 15442 22460
rect 18233 22457 18245 22460
rect 18279 22488 18291 22491
rect 18690 22488 18696 22500
rect 18279 22460 18696 22488
rect 18279 22457 18291 22460
rect 18233 22451 18291 22457
rect 18690 22448 18696 22460
rect 18748 22448 18754 22500
rect 18874 22448 18880 22500
rect 18932 22448 18938 22500
rect 7484 22392 10732 22420
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 10836 22392 10977 22420
rect 10836 22380 10842 22392
rect 10965 22389 10977 22392
rect 11011 22389 11023 22423
rect 10965 22383 11023 22389
rect 11698 22380 11704 22432
rect 11756 22380 11762 22432
rect 12526 22380 12532 22432
rect 12584 22420 12590 22432
rect 12621 22423 12679 22429
rect 12621 22420 12633 22423
rect 12584 22392 12633 22420
rect 12584 22380 12590 22392
rect 12621 22389 12633 22392
rect 12667 22389 12679 22423
rect 12621 22383 12679 22389
rect 12894 22380 12900 22432
rect 12952 22420 12958 22432
rect 19058 22420 19064 22432
rect 12952 22392 19064 22420
rect 12952 22380 12958 22392
rect 19058 22380 19064 22392
rect 19116 22380 19122 22432
rect 20530 22380 20536 22432
rect 20588 22380 20594 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 23569 22423 23627 22429
rect 23569 22389 23581 22423
rect 23615 22420 23627 22423
rect 24394 22420 24400 22432
rect 23615 22392 24400 22420
rect 23615 22389 23627 22392
rect 23569 22383 23627 22389
rect 24394 22380 24400 22392
rect 24452 22380 24458 22432
rect 26694 22380 26700 22432
rect 26752 22420 26758 22432
rect 27065 22423 27123 22429
rect 27065 22420 27077 22423
rect 26752 22392 27077 22420
rect 26752 22380 26758 22392
rect 27065 22389 27077 22392
rect 27111 22389 27123 22423
rect 27065 22383 27123 22389
rect 1104 22330 29716 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 29716 22330
rect 1104 22256 29716 22278
rect 3050 22176 3056 22228
rect 3108 22216 3114 22228
rect 4249 22219 4307 22225
rect 4249 22216 4261 22219
rect 3108 22188 4261 22216
rect 3108 22176 3114 22188
rect 4249 22185 4261 22188
rect 4295 22185 4307 22219
rect 4249 22179 4307 22185
rect 4433 22219 4491 22225
rect 4433 22185 4445 22219
rect 4479 22216 4491 22219
rect 4614 22216 4620 22228
rect 4479 22188 4620 22216
rect 4479 22185 4491 22188
rect 4433 22179 4491 22185
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 5258 22176 5264 22228
rect 5316 22216 5322 22228
rect 5316 22188 12664 22216
rect 5316 22176 5322 22188
rect 2958 22108 2964 22160
rect 3016 22148 3022 22160
rect 6546 22148 6552 22160
rect 3016 22120 6552 22148
rect 3016 22108 3022 22120
rect 6546 22108 6552 22120
rect 6604 22108 6610 22160
rect 6656 22120 7052 22148
rect 3881 22083 3939 22089
rect 3881 22049 3893 22083
rect 3927 22080 3939 22083
rect 4062 22080 4068 22092
rect 3927 22052 4068 22080
rect 3927 22049 3939 22052
rect 3881 22043 3939 22049
rect 4062 22040 4068 22052
rect 4120 22040 4126 22092
rect 6656 22080 6684 22120
rect 6380 22052 6684 22080
rect 6380 22021 6408 22052
rect 6822 22040 6828 22092
rect 6880 22040 6886 22092
rect 7024 22080 7052 22120
rect 7190 22108 7196 22160
rect 7248 22148 7254 22160
rect 7248 22120 7788 22148
rect 7248 22108 7254 22120
rect 7466 22080 7472 22092
rect 7024 22052 7472 22080
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 7650 22040 7656 22092
rect 7708 22040 7714 22092
rect 7760 22089 7788 22120
rect 8588 22120 9260 22148
rect 7745 22083 7803 22089
rect 7745 22049 7757 22083
rect 7791 22049 7803 22083
rect 8202 22080 8208 22092
rect 7745 22043 7803 22049
rect 7852 22052 8208 22080
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 22012 3847 22015
rect 6181 22015 6239 22021
rect 3835 21984 4108 22012
rect 3835 21981 3847 21984
rect 3789 21975 3847 21981
rect 4080 21956 4108 21984
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6181 21975 6239 21981
rect 6365 22015 6423 22021
rect 6365 21981 6377 22015
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 21981 6515 22015
rect 6457 21975 6515 21981
rect 6605 22015 6663 22021
rect 6605 21981 6617 22015
rect 6651 22012 6663 22015
rect 6651 21981 6684 22012
rect 6605 21975 6684 21981
rect 4062 21904 4068 21956
rect 4120 21904 4126 21956
rect 4617 21947 4675 21953
rect 4617 21944 4629 21947
rect 4264 21916 4629 21944
rect 3878 21836 3884 21888
rect 3936 21876 3942 21888
rect 4264 21876 4292 21916
rect 4617 21913 4629 21916
rect 4663 21944 4675 21947
rect 5350 21944 5356 21956
rect 4663 21916 5356 21944
rect 4663 21913 4675 21916
rect 4617 21907 4675 21913
rect 5350 21904 5356 21916
rect 5408 21904 5414 21956
rect 3936 21848 4292 21876
rect 4417 21879 4475 21885
rect 3936 21836 3942 21848
rect 4417 21845 4429 21879
rect 4463 21876 4475 21879
rect 4706 21876 4712 21888
rect 4463 21848 4712 21876
rect 4463 21845 4475 21848
rect 4417 21839 4475 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 6196 21876 6224 21975
rect 6273 21947 6331 21953
rect 6273 21913 6285 21947
rect 6319 21944 6331 21947
rect 6472 21944 6500 21975
rect 6319 21916 6500 21944
rect 6319 21913 6331 21916
rect 6273 21907 6331 21913
rect 6546 21876 6552 21888
rect 6196 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 6656 21876 6684 21975
rect 6730 21972 6736 22024
rect 6788 21972 6794 22024
rect 6840 22012 6868 22040
rect 6922 22015 6980 22021
rect 6922 22012 6934 22015
rect 6840 21984 6934 22012
rect 6922 21981 6934 21984
rect 6968 21981 6980 22015
rect 6922 21975 6980 21981
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 7561 22015 7619 22021
rect 7561 21981 7573 22015
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 6822 21904 6828 21956
rect 6880 21904 6886 21956
rect 7282 21944 7288 21956
rect 7024 21916 7288 21944
rect 7024 21876 7052 21916
rect 7282 21904 7288 21916
rect 7340 21904 7346 21956
rect 7576 21944 7604 21975
rect 7852 21944 7880 22052
rect 8202 22040 8208 22052
rect 8260 22040 8266 22092
rect 8478 22040 8484 22092
rect 8536 22080 8542 22092
rect 8588 22080 8616 22120
rect 8536 22052 8616 22080
rect 8536 22040 8542 22052
rect 8662 22040 8668 22092
rect 8720 22080 8726 22092
rect 9232 22089 9260 22120
rect 9646 22120 10180 22148
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 8720 22052 9076 22080
rect 9195 22052 9229 22080
rect 8720 22040 8726 22052
rect 7929 22015 7987 22021
rect 7929 21981 7941 22015
rect 7975 22012 7987 22015
rect 7975 21984 8064 22012
rect 7975 21981 7987 21984
rect 7929 21975 7987 21981
rect 7576 21916 7880 21944
rect 6656 21848 7052 21876
rect 7098 21836 7104 21888
rect 7156 21836 7162 21888
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 8036 21876 8064 21984
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 8573 22015 8631 22021
rect 8352 21984 8524 22012
rect 8352 21972 8358 21984
rect 8113 21947 8171 21953
rect 8113 21913 8125 21947
rect 8159 21944 8171 21947
rect 8205 21947 8263 21953
rect 8205 21944 8217 21947
rect 8159 21916 8217 21944
rect 8159 21913 8171 21916
rect 8113 21907 8171 21913
rect 8205 21913 8217 21916
rect 8251 21913 8263 21947
rect 8205 21907 8263 21913
rect 8386 21904 8392 21956
rect 8444 21904 8450 21956
rect 8496 21944 8524 21984
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8619 21984 8953 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 9048 22012 9076 22052
rect 9217 22049 9229 22052
rect 9263 22049 9275 22083
rect 9217 22043 9275 22049
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9646 22080 9674 22120
rect 9364 22052 9674 22080
rect 9364 22040 9370 22052
rect 9766 22040 9772 22092
rect 9824 22080 9830 22092
rect 9824 22052 10088 22080
rect 9824 22040 9830 22052
rect 9122 22012 9128 22024
rect 9048 21984 9128 22012
rect 8941 21975 8999 21981
rect 9122 21972 9128 21984
rect 9180 21972 9186 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 9232 21984 9505 22012
rect 9232 21944 9260 21984
rect 9493 21981 9505 21984
rect 9539 22012 9551 22015
rect 9539 21984 9904 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 8496 21916 9260 21944
rect 9398 21904 9404 21956
rect 9456 21944 9462 21956
rect 9456 21916 9812 21944
rect 9456 21904 9462 21916
rect 7984 21848 8064 21876
rect 7984 21836 7990 21848
rect 9582 21836 9588 21888
rect 9640 21876 9646 21888
rect 9784 21885 9812 21916
rect 9677 21879 9735 21885
rect 9677 21876 9689 21879
rect 9640 21848 9689 21876
rect 9640 21836 9646 21848
rect 9677 21845 9689 21848
rect 9723 21845 9735 21879
rect 9677 21839 9735 21845
rect 9769 21879 9827 21885
rect 9769 21845 9781 21879
rect 9815 21845 9827 21879
rect 9876 21876 9904 21984
rect 9950 21972 9956 22024
rect 10008 21972 10014 22024
rect 10060 22021 10088 22052
rect 10152 22021 10180 22120
rect 10226 22108 10232 22160
rect 10284 22148 10290 22160
rect 11333 22151 11391 22157
rect 11333 22148 11345 22151
rect 10284 22120 11345 22148
rect 10284 22108 10290 22120
rect 11333 22117 11345 22120
rect 11379 22117 11391 22151
rect 11333 22111 11391 22117
rect 11698 22108 11704 22160
rect 11756 22148 11762 22160
rect 12636 22148 12664 22188
rect 12710 22176 12716 22228
rect 12768 22216 12774 22228
rect 14829 22219 14887 22225
rect 12768 22188 14780 22216
rect 12768 22176 12774 22188
rect 12894 22148 12900 22160
rect 11756 22120 12480 22148
rect 12636 22120 12900 22148
rect 11756 22108 11762 22120
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 11517 22083 11575 22089
rect 10560 22052 10824 22080
rect 10560 22040 10566 22052
rect 10045 22015 10103 22021
rect 10045 21981 10057 22015
rect 10091 21981 10103 22015
rect 10045 21975 10103 21981
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10318 21972 10324 22024
rect 10376 21972 10382 22024
rect 10594 21972 10600 22024
rect 10652 22021 10658 22024
rect 10796 22021 10824 22052
rect 11164 22052 11468 22080
rect 10652 22015 10701 22021
rect 10652 21981 10655 22015
rect 10689 21981 10701 22015
rect 10652 21975 10701 21981
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 10652 21972 10658 21975
rect 10962 21972 10968 22024
rect 11020 22012 11026 22024
rect 11164 22021 11192 22052
rect 11056 22015 11114 22021
rect 11056 22012 11068 22015
rect 11020 21984 11068 22012
rect 11020 21972 11026 21984
rect 11056 21981 11068 21984
rect 11102 21981 11114 22015
rect 11056 21975 11114 21981
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 11238 21972 11244 22024
rect 11296 21972 11302 22024
rect 11440 22012 11468 22052
rect 11517 22049 11529 22083
rect 11563 22080 11575 22083
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 11563 22052 12357 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12452 22080 12480 22120
rect 12894 22108 12900 22120
rect 12952 22108 12958 22160
rect 13538 22108 13544 22160
rect 13596 22108 13602 22160
rect 14274 22108 14280 22160
rect 14332 22108 14338 22160
rect 14752 22148 14780 22188
rect 14829 22185 14841 22219
rect 14875 22216 14887 22219
rect 15194 22216 15200 22228
rect 14875 22188 15200 22216
rect 14875 22185 14887 22188
rect 14829 22179 14887 22185
rect 15194 22176 15200 22188
rect 15252 22176 15258 22228
rect 16945 22219 17003 22225
rect 16945 22185 16957 22219
rect 16991 22216 17003 22219
rect 17310 22216 17316 22228
rect 16991 22188 17316 22216
rect 16991 22185 17003 22188
rect 16945 22179 17003 22185
rect 17310 22176 17316 22188
rect 17368 22176 17374 22228
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20257 22219 20315 22225
rect 20257 22216 20269 22219
rect 20036 22188 20269 22216
rect 20036 22176 20042 22188
rect 20257 22185 20269 22188
rect 20303 22185 20315 22219
rect 20257 22179 20315 22185
rect 20530 22176 20536 22228
rect 20588 22216 20594 22228
rect 21158 22219 21216 22225
rect 21158 22216 21170 22219
rect 20588 22188 21170 22216
rect 20588 22176 20594 22188
rect 21158 22185 21170 22188
rect 21204 22185 21216 22219
rect 23842 22216 23848 22228
rect 21158 22179 21216 22185
rect 23308 22188 23848 22216
rect 20714 22148 20720 22160
rect 14752 22120 20720 22148
rect 12452 22052 13124 22080
rect 12345 22043 12403 22049
rect 11606 22012 11612 22024
rect 11440 21984 11612 22012
rect 11606 21972 11612 21984
rect 11664 21972 11670 22024
rect 11788 22015 11846 22021
rect 11788 21981 11800 22015
rect 11834 22012 11846 22015
rect 12066 22012 12072 22024
rect 11834 21984 12072 22012
rect 11834 21981 11846 21984
rect 11788 21975 11846 21981
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12160 22015 12218 22021
rect 12160 21981 12172 22015
rect 12206 21981 12218 22015
rect 12160 21975 12218 21981
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 22012 12311 22015
rect 12526 22012 12532 22024
rect 12584 22021 12590 22024
rect 13096 22021 13124 22052
rect 13354 22040 13360 22092
rect 13412 22040 13418 22092
rect 12584 22015 12617 22021
rect 12299 21984 12532 22012
rect 12299 21981 12311 21984
rect 12253 21975 12311 21981
rect 10873 21947 10931 21953
rect 10873 21913 10885 21947
rect 10919 21944 10931 21947
rect 11422 21944 11428 21956
rect 10919 21916 11428 21944
rect 10919 21913 10931 21916
rect 10873 21907 10931 21913
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 11882 21904 11888 21956
rect 11940 21904 11946 21956
rect 11974 21904 11980 21956
rect 12032 21904 12038 21956
rect 12176 21944 12204 21975
rect 12526 21972 12532 21984
rect 12605 21981 12617 22015
rect 12584 21975 12617 21981
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 21981 12771 22015
rect 12713 21975 12771 21981
rect 13081 22015 13139 22021
rect 13081 21981 13093 22015
rect 13127 21981 13139 22015
rect 13081 21975 13139 21981
rect 12584 21972 12590 21975
rect 12434 21944 12440 21956
rect 12176 21916 12440 21944
rect 12434 21904 12440 21916
rect 12492 21904 12498 21956
rect 12728 21944 12756 21975
rect 13170 21972 13176 22024
rect 13228 21972 13234 22024
rect 13262 21972 13268 22024
rect 13320 22012 13326 22024
rect 13556 22021 13584 22108
rect 14553 22083 14611 22089
rect 14553 22049 14565 22083
rect 14599 22080 14611 22083
rect 14826 22080 14832 22092
rect 14599 22052 14832 22080
rect 14599 22049 14611 22052
rect 14553 22043 14611 22049
rect 14826 22040 14832 22052
rect 14884 22080 14890 22092
rect 14884 22052 19288 22080
rect 14884 22040 14890 22052
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13320 21984 13461 22012
rect 13320 21972 13326 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 21981 13599 22015
rect 13541 21975 13599 21981
rect 13722 21972 13728 22024
rect 13780 21972 13786 22024
rect 14182 21972 14188 22024
rect 14240 21972 14246 22024
rect 14458 21972 14464 22024
rect 14516 22012 14522 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14516 21984 14657 22012
rect 14516 21972 14522 21984
rect 14645 21981 14657 21984
rect 14691 21981 14703 22015
rect 14645 21975 14703 21981
rect 13633 21947 13691 21953
rect 13633 21944 13645 21947
rect 12728 21916 13645 21944
rect 10318 21876 10324 21888
rect 9876 21848 10324 21876
rect 9769 21839 9827 21845
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 10505 21879 10563 21885
rect 10505 21845 10517 21879
rect 10551 21876 10563 21879
rect 11238 21876 11244 21888
rect 10551 21848 11244 21876
rect 10551 21845 10563 21848
rect 10505 21839 10563 21845
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 11514 21836 11520 21888
rect 11572 21836 11578 21888
rect 11606 21836 11612 21888
rect 11664 21836 11670 21888
rect 11698 21836 11704 21888
rect 11756 21876 11762 21888
rect 12728 21876 12756 21916
rect 13633 21913 13645 21916
rect 13679 21913 13691 21947
rect 14660 21944 14688 21975
rect 14734 21972 14740 22024
rect 14792 22012 14798 22024
rect 14918 22012 14924 22024
rect 14792 21984 14924 22012
rect 14792 21972 14798 21984
rect 14918 21972 14924 21984
rect 14976 21972 14982 22024
rect 15197 22015 15255 22021
rect 15197 21981 15209 22015
rect 15243 22012 15255 22015
rect 15378 22012 15384 22024
rect 15243 21984 15384 22012
rect 15243 21981 15255 21984
rect 15197 21975 15255 21981
rect 15378 21972 15384 21984
rect 15436 22012 15442 22024
rect 15654 22012 15660 22024
rect 15436 21984 15660 22012
rect 15436 21972 15442 21984
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 16853 22015 16911 22021
rect 16853 22012 16865 22015
rect 16816 21984 16865 22012
rect 16816 21972 16822 21984
rect 16853 21981 16865 21984
rect 16899 22012 16911 22015
rect 17126 22012 17132 22024
rect 16899 21984 17132 22012
rect 16899 21981 16911 21984
rect 16853 21975 16911 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 14826 21944 14832 21956
rect 14660 21916 14832 21944
rect 13633 21907 13691 21913
rect 14826 21904 14832 21916
rect 14884 21904 14890 21956
rect 19150 21944 19156 21956
rect 14936 21916 19156 21944
rect 11756 21848 12756 21876
rect 11756 21836 11762 21848
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14936 21876 14964 21916
rect 19150 21904 19156 21916
rect 19208 21904 19214 21956
rect 13964 21848 14964 21876
rect 13964 21836 13970 21848
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 17218 21836 17224 21888
rect 17276 21876 17282 21888
rect 17402 21876 17408 21888
rect 17276 21848 17408 21876
rect 17276 21836 17282 21848
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 19260 21876 19288 22052
rect 19518 22040 19524 22092
rect 19576 22040 19582 22092
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19392 21984 19441 22012
rect 19392 21972 19398 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19334 21876 19340 21888
rect 19260 21848 19340 21876
rect 19334 21836 19340 21848
rect 19392 21836 19398 21888
rect 19444 21876 19472 21975
rect 19702 21972 19708 22024
rect 19760 21972 19766 22024
rect 19812 21944 19840 22120
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 23308 22157 23336 22188
rect 23842 22176 23848 22188
rect 23900 22176 23906 22228
rect 24857 22219 24915 22225
rect 24857 22185 24869 22219
rect 24903 22216 24915 22219
rect 25298 22219 25356 22225
rect 25298 22216 25310 22219
rect 24903 22188 25310 22216
rect 24903 22185 24915 22188
rect 24857 22179 24915 22185
rect 25298 22185 25310 22188
rect 25344 22185 25356 22219
rect 25298 22179 25356 22185
rect 27154 22176 27160 22228
rect 27212 22216 27218 22228
rect 27433 22219 27491 22225
rect 27433 22216 27445 22219
rect 27212 22188 27445 22216
rect 27212 22176 27218 22188
rect 27433 22185 27445 22188
rect 27479 22185 27491 22219
rect 27433 22179 27491 22185
rect 23293 22151 23351 22157
rect 23293 22117 23305 22151
rect 23339 22117 23351 22151
rect 23293 22111 23351 22117
rect 23382 22108 23388 22160
rect 23440 22148 23446 22160
rect 23440 22120 24624 22148
rect 23440 22108 23446 22120
rect 20901 22083 20959 22089
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 21726 22080 21732 22092
rect 20947 22052 21732 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 21726 22040 21732 22052
rect 21784 22040 21790 22092
rect 21818 22040 21824 22092
rect 21876 22080 21882 22092
rect 22554 22080 22560 22092
rect 21876 22052 22560 22080
rect 21876 22040 21882 22052
rect 22554 22040 22560 22052
rect 22612 22080 22618 22092
rect 22612 22052 22968 22080
rect 22612 22040 22618 22052
rect 20070 21972 20076 22024
rect 20128 22012 20134 22024
rect 20254 22012 20260 22024
rect 20128 21984 20260 22012
rect 20128 21972 20134 21984
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 22940 22021 22968 22052
rect 24486 22040 24492 22092
rect 24544 22040 24550 22092
rect 24596 22080 24624 22120
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24596 22052 25053 22080
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 26050 22040 26056 22092
rect 26108 22080 26114 22092
rect 26108 22052 27292 22080
rect 26108 22040 26114 22052
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 19886 21944 19892 21956
rect 19812 21916 19892 21944
rect 19886 21904 19892 21916
rect 19944 21904 19950 21956
rect 19981 21947 20039 21953
rect 19981 21913 19993 21947
rect 20027 21944 20039 21947
rect 20162 21944 20168 21956
rect 20027 21916 20168 21944
rect 20027 21913 20039 21916
rect 19981 21907 20039 21913
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 22833 21947 22891 21953
rect 22833 21944 22845 21947
rect 22402 21916 22845 21944
rect 22833 21913 22845 21916
rect 22879 21913 22891 21947
rect 22833 21907 22891 21913
rect 23566 21904 23572 21956
rect 23624 21904 23630 21956
rect 20622 21876 20628 21888
rect 19444 21848 20628 21876
rect 20622 21836 20628 21848
rect 20680 21836 20686 21888
rect 22649 21879 22707 21885
rect 22649 21845 22661 21879
rect 22695 21876 22707 21879
rect 22922 21876 22928 21888
rect 22695 21848 22928 21876
rect 22695 21845 22707 21848
rect 22649 21839 22707 21845
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 23106 21836 23112 21888
rect 23164 21836 23170 21888
rect 24596 21876 24624 21975
rect 26602 21972 26608 22024
rect 26660 22012 26666 22024
rect 27264 22021 27292 22052
rect 28902 22040 28908 22092
rect 28960 22040 28966 22092
rect 27065 22015 27123 22021
rect 27065 22012 27077 22015
rect 26660 21984 27077 22012
rect 26660 21972 26666 21984
rect 27065 21981 27077 21984
rect 27111 21981 27123 22015
rect 27065 21975 27123 21981
rect 27249 22015 27307 22021
rect 27249 21981 27261 22015
rect 27295 21981 27307 22015
rect 27249 21975 27307 21981
rect 28994 21972 29000 22024
rect 29052 21972 29058 22024
rect 29270 21972 29276 22024
rect 29328 21972 29334 22024
rect 26694 21944 26700 21956
rect 26542 21916 26700 21944
rect 26694 21904 26700 21916
rect 26752 21904 26758 21956
rect 26881 21947 26939 21953
rect 26881 21913 26893 21947
rect 26927 21913 26939 21947
rect 26881 21907 26939 21913
rect 26789 21879 26847 21885
rect 26789 21876 26801 21879
rect 24596 21848 26801 21876
rect 26789 21845 26801 21848
rect 26835 21876 26847 21879
rect 26896 21876 26924 21907
rect 27062 21876 27068 21888
rect 26835 21848 27068 21876
rect 26835 21845 26847 21848
rect 26789 21839 26847 21845
rect 27062 21836 27068 21848
rect 27120 21836 27126 21888
rect 27154 21836 27160 21888
rect 27212 21836 27218 21888
rect 29178 21836 29184 21888
rect 29236 21836 29242 21888
rect 1104 21786 29716 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 29716 21786
rect 1104 21712 29716 21734
rect 6638 21672 6644 21684
rect 5828 21644 6644 21672
rect 3878 21564 3884 21616
rect 3936 21564 3942 21616
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 900 21508 1501 21536
rect 900 21496 906 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 2774 21496 2780 21548
rect 2832 21536 2838 21548
rect 2869 21539 2927 21545
rect 2869 21536 2881 21539
rect 2832 21508 2881 21536
rect 2832 21496 2838 21508
rect 2869 21505 2881 21508
rect 2915 21505 2927 21539
rect 2869 21499 2927 21505
rect 5534 21496 5540 21548
rect 5592 21536 5598 21548
rect 5721 21539 5779 21545
rect 5721 21536 5733 21539
rect 5592 21508 5733 21536
rect 5592 21496 5598 21508
rect 5721 21505 5733 21508
rect 5767 21536 5779 21539
rect 5828 21536 5856 21644
rect 6638 21632 6644 21644
rect 6696 21632 6702 21684
rect 7926 21672 7932 21684
rect 7484 21644 7932 21672
rect 5994 21564 6000 21616
rect 6052 21604 6058 21616
rect 6733 21607 6791 21613
rect 6733 21604 6745 21607
rect 6052 21576 6745 21604
rect 6052 21564 6058 21576
rect 6733 21573 6745 21576
rect 6779 21573 6791 21607
rect 6733 21567 6791 21573
rect 5767 21508 5856 21536
rect 5905 21539 5963 21545
rect 5767 21505 5779 21508
rect 5721 21499 5779 21505
rect 5905 21505 5917 21539
rect 5951 21536 5963 21539
rect 6454 21536 6460 21548
rect 5951 21508 6460 21536
rect 5951 21505 5963 21508
rect 5905 21499 5963 21505
rect 6454 21496 6460 21508
rect 6512 21536 6518 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 6638 21496 6644 21548
rect 6696 21496 6702 21548
rect 7484 21545 7512 21644
rect 7926 21632 7932 21644
rect 7984 21632 7990 21684
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 8386 21672 8392 21684
rect 8067 21644 8392 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 8386 21632 8392 21644
rect 8444 21632 8450 21684
rect 8573 21675 8631 21681
rect 8573 21641 8585 21675
rect 8619 21641 8631 21675
rect 8573 21635 8631 21641
rect 9493 21675 9551 21681
rect 9493 21641 9505 21675
rect 9539 21672 9551 21675
rect 10226 21672 10232 21684
rect 9539 21644 10232 21672
rect 9539 21641 9551 21644
rect 9493 21635 9551 21641
rect 7745 21607 7803 21613
rect 7745 21573 7757 21607
rect 7791 21604 7803 21607
rect 8478 21604 8484 21616
rect 7791 21576 8484 21604
rect 7791 21573 7803 21576
rect 7745 21567 7803 21573
rect 6917 21539 6975 21545
rect 6917 21505 6929 21539
rect 6963 21536 6975 21539
rect 7469 21539 7527 21545
rect 7469 21536 7481 21539
rect 6963 21508 7481 21536
rect 6963 21505 6975 21508
rect 6917 21499 6975 21505
rect 7469 21505 7481 21508
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 7653 21539 7711 21545
rect 7653 21505 7665 21539
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 3142 21428 3148 21480
rect 3200 21428 3206 21480
rect 4614 21428 4620 21480
rect 4672 21468 4678 21480
rect 4893 21471 4951 21477
rect 4893 21468 4905 21471
rect 4672 21440 4905 21468
rect 4672 21428 4678 21440
rect 4893 21437 4905 21440
rect 4939 21468 4951 21471
rect 6932 21468 6960 21499
rect 4939 21440 6960 21468
rect 4939 21437 4951 21440
rect 4893 21431 4951 21437
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 7668 21468 7696 21499
rect 7248 21440 7696 21468
rect 7248 21428 7254 21440
rect 1673 21403 1731 21409
rect 1673 21369 1685 21403
rect 1719 21400 1731 21403
rect 1762 21400 1768 21412
rect 1719 21372 1768 21400
rect 1719 21369 1731 21372
rect 1673 21363 1731 21369
rect 1762 21360 1768 21372
rect 1820 21360 1826 21412
rect 5905 21403 5963 21409
rect 5905 21369 5917 21403
rect 5951 21400 5963 21403
rect 6546 21400 6552 21412
rect 5951 21372 6552 21400
rect 5951 21369 5963 21372
rect 5905 21363 5963 21369
rect 6546 21360 6552 21372
rect 6604 21360 6610 21412
rect 6638 21360 6644 21412
rect 6696 21400 6702 21412
rect 7760 21400 7788 21567
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 8588 21604 8616 21635
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 11606 21672 11612 21684
rect 10652 21644 11612 21672
rect 10652 21632 10658 21644
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 15286 21632 15292 21684
rect 15344 21672 15350 21684
rect 15562 21672 15568 21684
rect 15344 21644 15568 21672
rect 15344 21632 15350 21644
rect 15562 21632 15568 21644
rect 15620 21672 15626 21684
rect 15620 21644 19012 21672
rect 15620 21632 15626 21644
rect 13173 21607 13231 21613
rect 8588 21576 11100 21604
rect 7837 21539 7895 21545
rect 7837 21505 7849 21539
rect 7883 21505 7895 21539
rect 7837 21499 7895 21505
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21505 8263 21539
rect 8205 21499 8263 21505
rect 6696 21372 7788 21400
rect 7852 21400 7880 21499
rect 8220 21468 8248 21499
rect 8386 21496 8392 21548
rect 8444 21496 8450 21548
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 8849 21539 8907 21545
rect 8849 21536 8861 21539
rect 8628 21508 8861 21536
rect 8628 21496 8634 21508
rect 8849 21505 8861 21508
rect 8895 21505 8907 21539
rect 8849 21499 8907 21505
rect 9398 21496 9404 21548
rect 9456 21496 9462 21548
rect 9582 21496 9588 21548
rect 9640 21496 9646 21548
rect 10594 21536 10600 21548
rect 9876 21508 10600 21536
rect 9876 21468 9904 21508
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 11072 21545 11100 21576
rect 13173 21573 13185 21607
rect 13219 21604 13231 21607
rect 13446 21604 13452 21616
rect 13219 21576 13452 21604
rect 13219 21573 13231 21576
rect 13173 21567 13231 21573
rect 13446 21564 13452 21576
rect 13504 21564 13510 21616
rect 14274 21564 14280 21616
rect 14332 21604 14338 21616
rect 14829 21607 14887 21613
rect 14829 21604 14841 21607
rect 14332 21576 14841 21604
rect 14332 21564 14338 21576
rect 14829 21573 14841 21576
rect 14875 21573 14887 21607
rect 16301 21607 16359 21613
rect 16301 21604 16313 21607
rect 14829 21567 14887 21573
rect 14936 21576 15332 21604
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21536 10747 21539
rect 11057 21539 11115 21545
rect 10735 21508 11008 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 8220 21440 9904 21468
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 10781 21471 10839 21477
rect 10781 21468 10793 21471
rect 10008 21440 10793 21468
rect 10008 21428 10014 21440
rect 10781 21437 10793 21440
rect 10827 21437 10839 21471
rect 10980 21468 11008 21508
rect 11057 21505 11069 21539
rect 11103 21505 11115 21539
rect 11057 21499 11115 21505
rect 11606 21496 11612 21548
rect 11664 21536 11670 21548
rect 11974 21536 11980 21548
rect 11664 21508 11980 21536
rect 11664 21496 11670 21508
rect 11974 21496 11980 21508
rect 12032 21496 12038 21548
rect 12986 21496 12992 21548
rect 13044 21496 13050 21548
rect 13081 21539 13139 21545
rect 13081 21505 13093 21539
rect 13127 21505 13139 21539
rect 13081 21499 13139 21505
rect 12526 21468 12532 21480
rect 10980 21440 12532 21468
rect 10781 21431 10839 21437
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 12618 21428 12624 21480
rect 12676 21468 12682 21480
rect 13096 21468 13124 21499
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 13320 21508 13369 21536
rect 13320 21496 13326 21508
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 14369 21539 14427 21545
rect 14369 21505 14381 21539
rect 14415 21505 14427 21539
rect 14369 21499 14427 21505
rect 13722 21468 13728 21480
rect 12676 21440 13728 21468
rect 12676 21428 12682 21440
rect 13722 21428 13728 21440
rect 13780 21428 13786 21480
rect 14384 21468 14412 21499
rect 14550 21496 14556 21548
rect 14608 21496 14614 21548
rect 14645 21539 14703 21545
rect 14645 21505 14657 21539
rect 14691 21536 14703 21539
rect 14734 21536 14740 21548
rect 14691 21508 14740 21536
rect 14691 21505 14703 21508
rect 14645 21499 14703 21505
rect 14734 21496 14740 21508
rect 14792 21496 14798 21548
rect 14936 21545 14964 21576
rect 14921 21539 14979 21545
rect 14921 21505 14933 21539
rect 14967 21505 14979 21539
rect 14921 21499 14979 21505
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 15194 21536 15200 21548
rect 15059 21508 15200 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 14936 21468 14964 21499
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15304 21545 15332 21576
rect 16132 21576 16313 21604
rect 15289 21539 15347 21545
rect 15289 21505 15301 21539
rect 15335 21536 15347 21539
rect 15470 21536 15476 21548
rect 15335 21508 15476 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 14384 21440 14964 21468
rect 15212 21468 15240 21496
rect 15381 21471 15439 21477
rect 15381 21468 15393 21471
rect 15212 21440 15393 21468
rect 15381 21437 15393 21440
rect 15427 21437 15439 21471
rect 15381 21431 15439 21437
rect 15562 21428 15568 21480
rect 15620 21428 15626 21480
rect 16132 21468 16160 21576
rect 16301 21573 16313 21576
rect 16347 21573 16359 21607
rect 16301 21567 16359 21573
rect 16390 21564 16396 21616
rect 16448 21604 16454 21616
rect 18984 21613 19012 21644
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 21140 21644 21189 21672
rect 21140 21632 21146 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 21913 21675 21971 21681
rect 21913 21641 21925 21675
rect 21959 21672 21971 21675
rect 22094 21672 22100 21684
rect 21959 21644 22100 21672
rect 21959 21641 21971 21644
rect 21913 21635 21971 21641
rect 22094 21632 22100 21644
rect 22152 21632 22158 21684
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 26234 21672 26240 21684
rect 24544 21644 26240 21672
rect 24544 21632 24550 21644
rect 26234 21632 26240 21644
rect 26292 21672 26298 21684
rect 26421 21675 26479 21681
rect 26421 21672 26433 21675
rect 26292 21644 26433 21672
rect 26292 21632 26298 21644
rect 26421 21641 26433 21644
rect 26467 21641 26479 21675
rect 26421 21635 26479 21641
rect 27154 21632 27160 21684
rect 27212 21672 27218 21684
rect 29273 21675 29331 21681
rect 29273 21672 29285 21675
rect 27212 21644 29285 21672
rect 27212 21632 27218 21644
rect 29273 21641 29285 21644
rect 29319 21641 29331 21675
rect 29273 21635 29331 21641
rect 16485 21607 16543 21613
rect 16485 21604 16497 21607
rect 16448 21576 16497 21604
rect 16448 21564 16454 21576
rect 16485 21573 16497 21576
rect 16531 21604 16543 21607
rect 17405 21607 17463 21613
rect 17405 21604 17417 21607
rect 16531 21576 17417 21604
rect 16531 21573 16543 21576
rect 16485 21567 16543 21573
rect 17405 21573 17417 21576
rect 17451 21573 17463 21607
rect 18969 21607 19027 21613
rect 17405 21567 17463 21573
rect 18524 21576 18920 21604
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21536 16267 21539
rect 16850 21536 16856 21548
rect 16255 21508 16856 21536
rect 16255 21505 16267 21508
rect 16209 21499 16267 21505
rect 16850 21496 16856 21508
rect 16908 21496 16914 21548
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21536 17003 21539
rect 16991 21508 17172 21536
rect 16991 21505 17003 21508
rect 16945 21499 17003 21505
rect 17144 21468 17172 21508
rect 17218 21496 17224 21548
rect 17276 21496 17282 21548
rect 17310 21496 17316 21548
rect 17368 21496 17374 21548
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21536 17555 21539
rect 17678 21536 17684 21548
rect 17543 21508 17684 21536
rect 17543 21505 17555 21508
rect 17497 21499 17555 21505
rect 17678 21496 17684 21508
rect 17736 21496 17742 21548
rect 18524 21545 18552 21576
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 18782 21496 18788 21548
rect 18840 21496 18846 21548
rect 18892 21536 18920 21576
rect 18969 21573 18981 21607
rect 19015 21573 19027 21607
rect 18969 21567 19027 21573
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 25409 21607 25467 21613
rect 21048 21576 21864 21604
rect 21048 21564 21054 21576
rect 21836 21548 21864 21576
rect 25409 21573 25421 21607
rect 25455 21604 25467 21607
rect 26326 21604 26332 21616
rect 25455 21576 26332 21604
rect 25455 21573 25467 21576
rect 25409 21567 25467 21573
rect 26326 21564 26332 21576
rect 26384 21604 26390 21616
rect 26384 21576 27568 21604
rect 26384 21564 26390 21576
rect 27540 21548 27568 21576
rect 28810 21564 28816 21616
rect 28868 21564 28874 21616
rect 19058 21536 19064 21548
rect 18892 21508 19064 21536
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 19518 21536 19524 21548
rect 19199 21508 19524 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 19518 21496 19524 21508
rect 19576 21496 19582 21548
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 20956 21508 21281 21536
rect 20956 21496 20962 21508
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 21818 21496 21824 21548
rect 21876 21496 21882 21548
rect 22922 21496 22928 21548
rect 22980 21496 22986 21548
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23198 21496 23204 21548
rect 23256 21496 23262 21548
rect 23345 21539 23403 21545
rect 23345 21505 23357 21539
rect 23391 21536 23403 21539
rect 23474 21536 23480 21548
rect 23391 21508 23480 21536
rect 23391 21505 23403 21508
rect 23345 21499 23403 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 24210 21536 24216 21548
rect 23716 21508 24216 21536
rect 23716 21496 23722 21508
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 25501 21539 25559 21545
rect 25501 21505 25513 21539
rect 25547 21505 25559 21539
rect 25501 21499 25559 21505
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21536 25927 21539
rect 26145 21539 26203 21545
rect 26145 21536 26157 21539
rect 25915 21508 26157 21536
rect 25915 21505 25927 21508
rect 25869 21499 25927 21505
rect 26145 21505 26157 21508
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 16132 21440 17172 21468
rect 17696 21468 17724 21496
rect 19978 21468 19984 21480
rect 17696 21440 19984 21468
rect 8757 21403 8815 21409
rect 8757 21400 8769 21403
rect 7852 21372 8769 21400
rect 6696 21360 6702 21372
rect 8757 21369 8769 21372
rect 8803 21400 8815 21403
rect 9122 21400 9128 21412
rect 8803 21372 9128 21400
rect 8803 21369 8815 21372
rect 8757 21363 8815 21369
rect 9122 21360 9128 21372
rect 9180 21360 9186 21412
rect 10965 21403 11023 21409
rect 10965 21369 10977 21403
rect 11011 21400 11023 21403
rect 11238 21400 11244 21412
rect 11011 21372 11244 21400
rect 11011 21369 11023 21372
rect 10965 21363 11023 21369
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 12544 21400 12572 21428
rect 13262 21400 13268 21412
rect 12544 21372 13268 21400
rect 13262 21360 13268 21372
rect 13320 21360 13326 21412
rect 15197 21403 15255 21409
rect 15197 21369 15209 21403
rect 15243 21400 15255 21403
rect 15580 21400 15608 21428
rect 15243 21372 15608 21400
rect 16485 21403 16543 21409
rect 15243 21369 15255 21372
rect 15197 21363 15255 21369
rect 16485 21369 16497 21403
rect 16531 21400 16543 21403
rect 17034 21400 17040 21412
rect 16531 21372 17040 21400
rect 16531 21369 16543 21372
rect 16485 21363 16543 21369
rect 17034 21360 17040 21372
rect 17092 21360 17098 21412
rect 17144 21400 17172 21440
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 18601 21403 18659 21409
rect 18601 21400 18613 21403
rect 17144 21372 18613 21400
rect 18601 21369 18613 21372
rect 18647 21400 18659 21403
rect 20806 21400 20812 21412
rect 18647 21372 20812 21400
rect 18647 21369 18659 21372
rect 18601 21363 18659 21369
rect 20806 21360 20812 21372
rect 20864 21360 20870 21412
rect 25516 21400 25544 21499
rect 25700 21468 25728 21499
rect 26234 21496 26240 21548
rect 26292 21496 26298 21548
rect 26418 21536 26424 21548
rect 26344 21508 26424 21536
rect 26344 21468 26372 21508
rect 26418 21496 26424 21508
rect 26476 21496 26482 21548
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21505 26663 21539
rect 26605 21499 26663 21505
rect 25700 21440 26372 21468
rect 26050 21400 26056 21412
rect 25516 21372 26056 21400
rect 26050 21360 26056 21372
rect 26108 21400 26114 21412
rect 26620 21400 26648 21499
rect 26970 21496 26976 21548
rect 27028 21496 27034 21548
rect 27522 21496 27528 21548
rect 27580 21496 27586 21548
rect 27433 21471 27491 21477
rect 27433 21437 27445 21471
rect 27479 21468 27491 21471
rect 27801 21471 27859 21477
rect 27801 21468 27813 21471
rect 27479 21440 27813 21468
rect 27479 21437 27491 21440
rect 27433 21431 27491 21437
rect 27801 21437 27813 21440
rect 27847 21437 27859 21471
rect 27801 21431 27859 21437
rect 26108 21372 26648 21400
rect 26108 21360 26114 21372
rect 27338 21360 27344 21412
rect 27396 21360 27402 21412
rect 6365 21335 6423 21341
rect 6365 21301 6377 21335
rect 6411 21332 6423 21335
rect 6822 21332 6828 21344
rect 6411 21304 6828 21332
rect 6411 21301 6423 21304
rect 6365 21295 6423 21301
rect 6822 21292 6828 21304
rect 6880 21292 6886 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 8205 21335 8263 21341
rect 8205 21332 8217 21335
rect 7432 21304 8217 21332
rect 7432 21292 7438 21304
rect 8205 21301 8217 21304
rect 8251 21301 8263 21335
rect 8205 21295 8263 21301
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 10502 21332 10508 21344
rect 8720 21304 10508 21332
rect 8720 21292 8726 21304
rect 10502 21292 10508 21304
rect 10560 21332 10566 21344
rect 10597 21335 10655 21341
rect 10597 21332 10609 21335
rect 10560 21304 10609 21332
rect 10560 21292 10566 21304
rect 10597 21301 10609 21304
rect 10643 21301 10655 21335
rect 10597 21295 10655 21301
rect 11057 21335 11115 21341
rect 11057 21301 11069 21335
rect 11103 21332 11115 21335
rect 11882 21332 11888 21344
rect 11103 21304 11888 21332
rect 11103 21301 11115 21304
rect 11057 21295 11115 21301
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 12805 21335 12863 21341
rect 12805 21301 12817 21335
rect 12851 21332 12863 21335
rect 13354 21332 13360 21344
rect 12851 21304 13360 21332
rect 12851 21301 12863 21304
rect 12805 21295 12863 21301
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14553 21335 14611 21341
rect 14553 21332 14565 21335
rect 14516 21304 14565 21332
rect 14516 21292 14522 21304
rect 14553 21301 14565 21304
rect 14599 21301 14611 21335
rect 14553 21295 14611 21301
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21332 15531 21335
rect 16298 21332 16304 21344
rect 15519 21304 16304 21332
rect 15519 21301 15531 21304
rect 15473 21295 15531 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 16669 21335 16727 21341
rect 16669 21332 16681 21335
rect 16632 21304 16681 21332
rect 16632 21292 16638 21304
rect 16669 21301 16681 21304
rect 16715 21301 16727 21335
rect 16669 21295 16727 21301
rect 17126 21292 17132 21344
rect 17184 21292 17190 21344
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 19058 21332 19064 21344
rect 17368 21304 19064 21332
rect 17368 21292 17374 21304
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 19337 21335 19395 21341
rect 19337 21301 19349 21335
rect 19383 21332 19395 21335
rect 19610 21332 19616 21344
rect 19383 21304 19616 21332
rect 19383 21301 19395 21304
rect 19337 21295 19395 21301
rect 19610 21292 19616 21304
rect 19668 21292 19674 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 23750 21332 23756 21344
rect 23523 21304 23756 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 25314 21292 25320 21344
rect 25372 21332 25378 21344
rect 25961 21335 26019 21341
rect 25961 21332 25973 21335
rect 25372 21304 25973 21332
rect 25372 21292 25378 21304
rect 25961 21301 25973 21304
rect 26007 21301 26019 21335
rect 25961 21295 26019 21301
rect 1104 21242 29716 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 29716 21242
rect 1104 21168 29716 21190
rect 3878 21088 3884 21140
rect 3936 21128 3942 21140
rect 4065 21131 4123 21137
rect 4065 21128 4077 21131
rect 3936 21100 4077 21128
rect 3936 21088 3942 21100
rect 4065 21097 4077 21100
rect 4111 21097 4123 21131
rect 4065 21091 4123 21097
rect 6270 21088 6276 21140
rect 6328 21128 6334 21140
rect 6730 21128 6736 21140
rect 6328 21100 6736 21128
rect 6328 21088 6334 21100
rect 6730 21088 6736 21100
rect 6788 21088 6794 21140
rect 7466 21088 7472 21140
rect 7524 21128 7530 21140
rect 8662 21128 8668 21140
rect 7524 21100 8668 21128
rect 7524 21088 7530 21100
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 9125 21131 9183 21137
rect 9125 21097 9137 21131
rect 9171 21128 9183 21131
rect 9306 21128 9312 21140
rect 9171 21100 9312 21128
rect 9171 21097 9183 21100
rect 9125 21091 9183 21097
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 9950 21088 9956 21140
rect 10008 21088 10014 21140
rect 12897 21131 12955 21137
rect 10060 21100 12112 21128
rect 6472 21032 9444 21060
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6178 20992 6184 21004
rect 5868 20964 6184 20992
rect 5868 20952 5874 20964
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6472 20936 6500 21032
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 8202 20992 8208 21004
rect 6972 20964 8208 20992
rect 6972 20952 6978 20964
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 4062 20884 4068 20936
rect 4120 20924 4126 20936
rect 6086 20933 6092 20936
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 4120 20896 4169 20924
rect 4120 20884 4126 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 6084 20924 6092 20933
rect 6047 20896 6092 20924
rect 4157 20887 4215 20893
rect 6084 20887 6092 20896
rect 6086 20884 6092 20887
rect 6144 20884 6150 20936
rect 6454 20924 6460 20936
rect 6415 20896 6460 20924
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 6546 20884 6552 20936
rect 6604 20884 6610 20936
rect 6822 20884 6828 20936
rect 6880 20884 6886 20936
rect 7282 20884 7288 20936
rect 7340 20924 7346 20936
rect 8386 20924 8392 20936
rect 7340 20896 8392 20924
rect 7340 20884 7346 20896
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 9214 20884 9220 20936
rect 9272 20884 9278 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 9416 20933 9444 21032
rect 9402 20927 9460 20933
rect 9402 20893 9414 20927
rect 9448 20924 9460 20927
rect 9490 20924 9496 20936
rect 9448 20896 9496 20924
rect 9448 20893 9460 20896
rect 9402 20887 9460 20893
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 9815 20927 9873 20933
rect 9815 20893 9827 20927
rect 9861 20924 9873 20927
rect 9950 20924 9956 20936
rect 9861 20896 9956 20924
rect 9861 20893 9873 20896
rect 9815 20887 9873 20893
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10060 20933 10088 21100
rect 11514 21020 11520 21072
rect 11572 21060 11578 21072
rect 11572 21032 12020 21060
rect 11572 21020 11578 21032
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20893 10103 20927
rect 10045 20887 10103 20893
rect 1394 20816 1400 20868
rect 1452 20856 1458 20868
rect 2774 20856 2780 20868
rect 1452 20828 2780 20856
rect 1452 20816 1458 20828
rect 2774 20816 2780 20828
rect 2832 20856 2838 20868
rect 3510 20856 3516 20868
rect 2832 20828 3516 20856
rect 2832 20816 2838 20828
rect 3510 20816 3516 20828
rect 3568 20856 3574 20868
rect 3568 20828 6040 20856
rect 3568 20816 3574 20828
rect 6012 20800 6040 20828
rect 6178 20816 6184 20868
rect 6236 20816 6242 20868
rect 6273 20859 6331 20865
rect 6273 20825 6285 20859
rect 6319 20856 6331 20859
rect 6362 20856 6368 20868
rect 6319 20828 6368 20856
rect 6319 20825 6331 20828
rect 6273 20819 6331 20825
rect 6362 20816 6368 20828
rect 6420 20816 6426 20868
rect 6914 20856 6920 20868
rect 6471 20828 6920 20856
rect 5902 20748 5908 20800
rect 5960 20748 5966 20800
rect 5994 20748 6000 20800
rect 6052 20788 6058 20800
rect 6471 20788 6499 20828
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 8665 20859 8723 20865
rect 8665 20825 8677 20859
rect 8711 20825 8723 20859
rect 8665 20819 8723 20825
rect 6052 20760 6499 20788
rect 6052 20748 6058 20760
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 6733 20791 6791 20797
rect 6733 20788 6745 20791
rect 6604 20760 6745 20788
rect 6604 20748 6610 20760
rect 6733 20757 6745 20760
rect 6779 20757 6791 20791
rect 8680 20788 8708 20819
rect 8938 20816 8944 20868
rect 8996 20856 9002 20868
rect 9585 20859 9643 20865
rect 9585 20856 9597 20859
rect 8996 20828 9597 20856
rect 8996 20816 9002 20828
rect 9585 20825 9597 20828
rect 9631 20825 9643 20859
rect 9585 20819 9643 20825
rect 9674 20816 9680 20868
rect 9732 20816 9738 20868
rect 10060 20788 10088 20887
rect 11882 20884 11888 20936
rect 11940 20884 11946 20936
rect 11992 20924 12020 21032
rect 12084 20992 12112 21100
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 12986 21128 12992 21140
rect 12943 21100 12992 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 17957 21131 18015 21137
rect 17957 21128 17969 21131
rect 15620 21100 17969 21128
rect 15620 21088 15626 21100
rect 17957 21097 17969 21100
rect 18003 21097 18015 21131
rect 20346 21128 20352 21140
rect 17957 21091 18015 21097
rect 18800 21100 20352 21128
rect 18800 21072 18828 21100
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 23198 21088 23204 21140
rect 23256 21088 23262 21140
rect 26418 21088 26424 21140
rect 26476 21128 26482 21140
rect 26789 21131 26847 21137
rect 26789 21128 26801 21131
rect 26476 21100 26801 21128
rect 26476 21088 26482 21100
rect 26789 21097 26801 21100
rect 26835 21097 26847 21131
rect 26789 21091 26847 21097
rect 12161 21063 12219 21069
rect 12161 21029 12173 21063
rect 12207 21060 12219 21063
rect 14366 21060 14372 21072
rect 12207 21032 14372 21060
rect 12207 21029 12219 21032
rect 12161 21023 12219 21029
rect 14366 21020 14372 21032
rect 14424 21020 14430 21072
rect 15470 21020 15476 21072
rect 15528 21060 15534 21072
rect 18782 21060 18788 21072
rect 15528 21032 18788 21060
rect 15528 21020 15534 21032
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 21082 21060 21088 21072
rect 19812 21032 21088 21060
rect 16482 20992 16488 21004
rect 12084 20964 16488 20992
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 17218 20952 17224 21004
rect 17276 20992 17282 21004
rect 17276 20964 18920 20992
rect 17276 20952 17282 20964
rect 12161 20927 12219 20933
rect 12161 20924 12173 20927
rect 11992 20896 12173 20924
rect 12161 20893 12173 20896
rect 12207 20893 12219 20927
rect 12161 20887 12219 20893
rect 12802 20884 12808 20936
rect 12860 20884 12866 20936
rect 16390 20884 16396 20936
rect 16448 20884 16454 20936
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 16853 20927 16911 20933
rect 16853 20924 16865 20927
rect 16632 20896 16865 20924
rect 16632 20884 16638 20896
rect 16853 20893 16865 20896
rect 16899 20893 16911 20927
rect 16853 20887 16911 20893
rect 17034 20884 17040 20936
rect 17092 20884 17098 20936
rect 17954 20884 17960 20936
rect 18012 20884 18018 20936
rect 18046 20884 18052 20936
rect 18104 20884 18110 20936
rect 10962 20816 10968 20868
rect 11020 20856 11026 20868
rect 11330 20856 11336 20868
rect 11020 20828 11336 20856
rect 11020 20816 11026 20828
rect 11330 20816 11336 20828
rect 11388 20856 11394 20868
rect 11790 20856 11796 20868
rect 11388 20828 11796 20856
rect 11388 20816 11394 20828
rect 11790 20816 11796 20828
rect 11848 20816 11854 20868
rect 16206 20816 16212 20868
rect 16264 20856 16270 20868
rect 16264 20828 16896 20856
rect 16264 20816 16270 20828
rect 16868 20800 16896 20828
rect 18230 20816 18236 20868
rect 18288 20816 18294 20868
rect 18892 20856 18920 20964
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19812 21001 19840 21032
rect 21082 21020 21088 21032
rect 21140 21020 21146 21072
rect 23566 21020 23572 21072
rect 23624 21020 23630 21072
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 19116 20964 19717 20992
rect 19116 20952 19122 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 19797 20995 19855 21001
rect 19797 20961 19809 20995
rect 19843 20961 19855 20995
rect 19797 20955 19855 20961
rect 20165 20995 20223 21001
rect 20165 20961 20177 20995
rect 20211 20992 20223 20995
rect 21453 20995 21511 21001
rect 20211 20964 21036 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 19518 20884 19524 20936
rect 19576 20924 19582 20936
rect 19613 20927 19671 20933
rect 19613 20924 19625 20927
rect 19576 20896 19625 20924
rect 19576 20884 19582 20896
rect 19613 20893 19625 20896
rect 19659 20893 19671 20927
rect 19613 20887 19671 20893
rect 19978 20884 19984 20936
rect 20036 20884 20042 20936
rect 20436 20927 20494 20933
rect 20436 20893 20448 20927
rect 20482 20924 20494 20927
rect 20482 20896 20760 20924
rect 20482 20893 20494 20896
rect 20436 20887 20494 20893
rect 20533 20859 20591 20865
rect 20533 20856 20545 20859
rect 18892 20828 20545 20856
rect 20533 20825 20545 20828
rect 20579 20825 20591 20859
rect 20533 20819 20591 20825
rect 20622 20816 20628 20868
rect 20680 20816 20686 20868
rect 8680 20760 10088 20788
rect 6733 20751 6791 20757
rect 11882 20748 11888 20800
rect 11940 20788 11946 20800
rect 11977 20791 12035 20797
rect 11977 20788 11989 20791
rect 11940 20760 11989 20788
rect 11940 20748 11946 20760
rect 11977 20757 11989 20760
rect 12023 20757 12035 20791
rect 11977 20751 12035 20757
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 13538 20788 13544 20800
rect 12492 20760 13544 20788
rect 12492 20748 12498 20760
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 16666 20748 16672 20800
rect 16724 20788 16730 20800
rect 16761 20791 16819 20797
rect 16761 20788 16773 20791
rect 16724 20760 16773 20788
rect 16724 20748 16730 20760
rect 16761 20757 16773 20760
rect 16807 20757 16819 20791
rect 16761 20751 16819 20757
rect 16850 20748 16856 20800
rect 16908 20748 16914 20800
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 17773 20791 17831 20797
rect 17773 20788 17785 20791
rect 17000 20760 17785 20788
rect 17000 20748 17006 20760
rect 17773 20757 17785 20760
rect 17819 20757 17831 20791
rect 17773 20751 17831 20757
rect 20254 20748 20260 20800
rect 20312 20748 20318 20800
rect 20732 20788 20760 20896
rect 20806 20884 20812 20936
rect 20864 20884 20870 20936
rect 21008 20933 21036 20964
rect 21453 20961 21465 20995
rect 21499 20992 21511 20995
rect 21726 20992 21732 21004
rect 21499 20964 21732 20992
rect 21499 20961 21511 20964
rect 21453 20955 21511 20961
rect 21726 20952 21732 20964
rect 21784 20992 21790 21004
rect 22094 20992 22100 21004
rect 21784 20964 22100 20992
rect 21784 20952 21790 20964
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 23934 20952 23940 21004
rect 23992 20952 23998 21004
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 26326 20992 26332 21004
rect 25087 20964 26332 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 26326 20952 26332 20964
rect 26384 20952 26390 21004
rect 26804 20992 26832 21091
rect 27338 21088 27344 21140
rect 27396 21128 27402 21140
rect 27433 21131 27491 21137
rect 27433 21128 27445 21131
rect 27396 21100 27445 21128
rect 27396 21088 27402 21100
rect 27433 21097 27445 21100
rect 27479 21097 27491 21131
rect 27433 21091 27491 21097
rect 28721 21131 28779 21137
rect 28721 21097 28733 21131
rect 28767 21128 28779 21131
rect 28810 21128 28816 21140
rect 28767 21100 28816 21128
rect 28767 21097 28779 21100
rect 28721 21091 28779 21097
rect 28810 21088 28816 21100
rect 28868 21088 28874 21140
rect 27157 20995 27215 21001
rect 27157 20992 27169 20995
rect 26804 20964 27169 20992
rect 27157 20961 27169 20964
rect 27203 20961 27215 20995
rect 27157 20955 27215 20961
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 20993 20927 21051 20933
rect 20993 20893 21005 20927
rect 21039 20893 21051 20927
rect 20993 20887 21051 20893
rect 20916 20856 20944 20887
rect 24394 20884 24400 20936
rect 24452 20884 24458 20936
rect 24486 20884 24492 20936
rect 24544 20924 24550 20936
rect 24673 20927 24731 20933
rect 24673 20924 24685 20927
rect 24544 20896 24685 20924
rect 24544 20884 24550 20896
rect 24673 20893 24685 20896
rect 24719 20893 24731 20927
rect 24673 20887 24731 20893
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20893 24823 20927
rect 24765 20887 24823 20893
rect 26973 20927 27031 20933
rect 26973 20893 26985 20927
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 21174 20856 21180 20868
rect 20916 20828 21180 20856
rect 21174 20816 21180 20828
rect 21232 20816 21238 20868
rect 21726 20816 21732 20868
rect 21784 20816 21790 20868
rect 22462 20816 22468 20868
rect 22520 20816 22526 20868
rect 23106 20816 23112 20868
rect 23164 20856 23170 20868
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 23164 20828 24593 20856
rect 23164 20816 23170 20828
rect 24581 20825 24593 20828
rect 24627 20825 24639 20859
rect 24581 20819 24639 20825
rect 20898 20788 20904 20800
rect 20732 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 20990 20748 20996 20800
rect 21048 20788 21054 20800
rect 21361 20791 21419 20797
rect 21361 20788 21373 20791
rect 21048 20760 21373 20788
rect 21048 20748 21054 20760
rect 21361 20757 21373 20760
rect 21407 20757 21419 20791
rect 21361 20751 21419 20757
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 24780 20788 24808 20887
rect 25314 20816 25320 20868
rect 25372 20816 25378 20868
rect 26326 20816 26332 20868
rect 26384 20816 26390 20868
rect 26988 20856 27016 20887
rect 27062 20884 27068 20936
rect 27120 20884 27126 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20893 27307 20927
rect 27249 20887 27307 20893
rect 28813 20927 28871 20933
rect 28813 20893 28825 20927
rect 28859 20924 28871 20927
rect 28994 20924 29000 20936
rect 28859 20896 29000 20924
rect 28859 20893 28871 20896
rect 28813 20887 28871 20893
rect 27154 20856 27160 20868
rect 26988 20828 27160 20856
rect 27154 20816 27160 20828
rect 27212 20816 27218 20868
rect 23532 20760 24808 20788
rect 23532 20748 23538 20760
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 24949 20791 25007 20797
rect 24949 20788 24961 20791
rect 24912 20760 24961 20788
rect 24912 20748 24918 20760
rect 24949 20757 24961 20760
rect 24995 20757 25007 20791
rect 24949 20751 25007 20757
rect 26050 20748 26056 20800
rect 26108 20788 26114 20800
rect 27264 20788 27292 20887
rect 28994 20884 29000 20896
rect 29052 20884 29058 20936
rect 29270 20884 29276 20936
rect 29328 20884 29334 20936
rect 26108 20760 27292 20788
rect 29181 20791 29239 20797
rect 26108 20748 26114 20760
rect 29181 20757 29193 20791
rect 29227 20788 29239 20791
rect 29822 20788 29828 20800
rect 29227 20760 29828 20788
rect 29227 20757 29239 20760
rect 29181 20751 29239 20757
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 1104 20698 29716 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 29716 20698
rect 1104 20624 29716 20646
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 6880 20556 8064 20584
rect 6880 20544 6886 20556
rect 4798 20476 4804 20528
rect 4856 20476 4862 20528
rect 6840 20516 6868 20544
rect 5920 20488 6868 20516
rect 3510 20408 3516 20460
rect 3568 20408 3574 20460
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 5920 20457 5948 20488
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 7745 20519 7803 20525
rect 7745 20516 7757 20519
rect 7156 20488 7757 20516
rect 7156 20476 7162 20488
rect 7745 20485 7757 20488
rect 7791 20485 7803 20519
rect 7745 20479 7803 20485
rect 5905 20451 5963 20457
rect 5905 20417 5917 20451
rect 5951 20417 5963 20451
rect 5905 20411 5963 20417
rect 6914 20408 6920 20460
rect 6972 20448 6978 20460
rect 8036 20457 8064 20556
rect 8404 20556 9260 20584
rect 7009 20451 7067 20457
rect 7009 20448 7021 20451
rect 6972 20420 7021 20448
rect 6972 20408 6978 20420
rect 7009 20417 7021 20420
rect 7055 20417 7067 20451
rect 8021 20451 8079 20457
rect 7009 20411 7067 20417
rect 7116 20420 7972 20448
rect 3786 20340 3792 20392
rect 3844 20340 3850 20392
rect 5534 20340 5540 20392
rect 5592 20340 5598 20392
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 7116 20380 7144 20420
rect 6236 20352 7144 20380
rect 6236 20340 6242 20352
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7248 20352 7849 20380
rect 7248 20340 7254 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7944 20380 7972 20420
rect 8021 20417 8033 20451
rect 8067 20417 8079 20451
rect 8021 20411 8079 20417
rect 8110 20408 8116 20460
rect 8168 20448 8174 20460
rect 8297 20451 8355 20457
rect 8297 20448 8309 20451
rect 8168 20420 8309 20448
rect 8168 20408 8174 20420
rect 8297 20417 8309 20420
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 8404 20380 8432 20556
rect 8570 20476 8576 20528
rect 8628 20516 8634 20528
rect 9033 20519 9091 20525
rect 9033 20516 9045 20519
rect 8628 20488 9045 20516
rect 8628 20476 8634 20488
rect 9033 20485 9045 20488
rect 9079 20485 9091 20519
rect 9232 20516 9260 20556
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 9401 20587 9459 20593
rect 9401 20584 9413 20587
rect 9364 20556 9413 20584
rect 9364 20544 9370 20556
rect 9401 20553 9413 20556
rect 9447 20553 9459 20587
rect 9401 20547 9459 20553
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 9548 20556 9812 20584
rect 9548 20544 9554 20556
rect 9674 20516 9680 20528
rect 9232 20488 9680 20516
rect 9033 20479 9091 20485
rect 8938 20457 8944 20460
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20417 8815 20451
rect 8757 20411 8815 20417
rect 8905 20451 8944 20457
rect 8905 20417 8917 20451
rect 8905 20411 8944 20417
rect 7944 20352 8432 20380
rect 8772 20380 8800 20411
rect 8938 20408 8944 20411
rect 8996 20408 9002 20460
rect 9122 20408 9128 20460
rect 9180 20408 9186 20460
rect 9214 20408 9220 20460
rect 9272 20457 9278 20460
rect 9508 20457 9536 20488
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 9272 20448 9280 20457
rect 9493 20451 9551 20457
rect 9272 20420 9317 20448
rect 9272 20411 9280 20420
rect 9493 20417 9505 20451
rect 9539 20417 9551 20451
rect 9493 20411 9551 20417
rect 9272 20408 9278 20411
rect 9784 20392 9812 20556
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 12989 20587 13047 20593
rect 10836 20556 12940 20584
rect 10836 20544 10842 20556
rect 9861 20519 9919 20525
rect 9861 20485 9873 20519
rect 9907 20516 9919 20519
rect 10042 20516 10048 20528
rect 9907 20488 10048 20516
rect 9907 20485 9919 20488
rect 9861 20479 9919 20485
rect 10042 20476 10048 20488
rect 10100 20516 10106 20528
rect 10686 20516 10692 20528
rect 10100 20488 10692 20516
rect 10100 20476 10106 20488
rect 10686 20476 10692 20488
rect 10744 20476 10750 20528
rect 11698 20516 11704 20528
rect 11256 20488 11704 20516
rect 10226 20448 10232 20460
rect 9876 20420 10232 20448
rect 9876 20392 9904 20420
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 9398 20380 9404 20392
rect 8772 20352 9404 20380
rect 7837 20343 7895 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9508 20352 9597 20380
rect 9508 20324 9536 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 9766 20380 9772 20392
rect 9723 20352 9772 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 9766 20340 9772 20352
rect 9824 20340 9830 20392
rect 9858 20340 9864 20392
rect 9916 20340 9922 20392
rect 11256 20380 11284 20488
rect 11698 20476 11704 20488
rect 11756 20476 11762 20528
rect 11793 20519 11851 20525
rect 11793 20485 11805 20519
rect 11839 20516 11851 20519
rect 12158 20516 12164 20528
rect 11839 20488 12164 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 12158 20476 12164 20488
rect 12216 20476 12222 20528
rect 12912 20516 12940 20556
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13449 20587 13507 20593
rect 13449 20584 13461 20587
rect 13035 20556 13461 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13449 20553 13461 20556
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14323 20556 14504 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 12912 20488 13492 20516
rect 11330 20408 11336 20460
rect 11388 20448 11394 20460
rect 11885 20451 11943 20457
rect 11388 20438 11744 20448
rect 11885 20438 11897 20451
rect 11388 20420 11897 20438
rect 11388 20408 11394 20420
rect 11716 20417 11897 20420
rect 11931 20417 11943 20451
rect 11716 20411 11943 20417
rect 11716 20410 11928 20411
rect 11974 20408 11980 20460
rect 12032 20408 12038 20460
rect 12342 20448 12348 20460
rect 12176 20420 12348 20448
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 11072 20352 11529 20380
rect 6012 20284 7788 20312
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 6012 20253 6040 20284
rect 5997 20247 6055 20253
rect 5997 20244 6009 20247
rect 5960 20216 6009 20244
rect 5960 20204 5966 20216
rect 5997 20213 6009 20216
rect 6043 20213 6055 20247
rect 5997 20207 6055 20213
rect 6181 20247 6239 20253
rect 6181 20213 6193 20247
rect 6227 20244 6239 20247
rect 6362 20244 6368 20256
rect 6227 20216 6368 20244
rect 6227 20213 6239 20216
rect 6181 20207 6239 20213
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 7760 20253 7788 20284
rect 7926 20272 7932 20324
rect 7984 20312 7990 20324
rect 8110 20312 8116 20324
rect 7984 20284 8116 20312
rect 7984 20272 7990 20284
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 8386 20272 8392 20324
rect 8444 20272 8450 20324
rect 9030 20272 9036 20324
rect 9088 20312 9094 20324
rect 9490 20312 9496 20324
rect 9088 20284 9496 20312
rect 9088 20272 9094 20284
rect 9490 20272 9496 20284
rect 9548 20272 9554 20324
rect 11072 20312 11100 20352
rect 11517 20349 11529 20352
rect 11563 20349 11575 20383
rect 11517 20343 11575 20349
rect 11609 20383 11667 20389
rect 11609 20349 11621 20383
rect 11655 20380 11667 20383
rect 12176 20380 12204 20420
rect 12342 20408 12348 20420
rect 12400 20448 12406 20460
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 12400 20420 12541 20448
rect 12400 20408 12406 20420
rect 12529 20417 12541 20420
rect 12575 20448 12587 20451
rect 12575 20420 13032 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 11655 20352 12204 20380
rect 12253 20383 12311 20389
rect 11655 20349 11667 20352
rect 11609 20343 11667 20349
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 12872 20383 12930 20389
rect 12872 20380 12884 20383
rect 12299 20352 12884 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 12872 20349 12884 20352
rect 12918 20349 12930 20383
rect 13004 20380 13032 20420
rect 13078 20408 13084 20460
rect 13136 20408 13142 20460
rect 13354 20408 13360 20460
rect 13412 20408 13418 20460
rect 13464 20457 13492 20488
rect 13814 20476 13820 20528
rect 13872 20476 13878 20528
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13688 20420 13737 20448
rect 13688 20408 13694 20420
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 13906 20408 13912 20460
rect 13964 20408 13970 20460
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 14476 20457 14504 20556
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 15105 20587 15163 20593
rect 14608 20556 14780 20584
rect 14608 20544 14614 20556
rect 14752 20525 14780 20556
rect 15105 20553 15117 20587
rect 15151 20584 15163 20587
rect 19061 20587 19119 20593
rect 15151 20556 16068 20584
rect 15151 20553 15163 20556
rect 15105 20547 15163 20553
rect 14737 20519 14795 20525
rect 14737 20485 14749 20519
rect 14783 20485 14795 20519
rect 14737 20479 14795 20485
rect 14829 20519 14887 20525
rect 14829 20485 14841 20519
rect 14875 20516 14887 20519
rect 15010 20516 15016 20528
rect 14875 20488 15016 20516
rect 14875 20485 14887 20488
rect 14829 20479 14887 20485
rect 15010 20476 15016 20488
rect 15068 20516 15074 20528
rect 16040 20525 16068 20556
rect 19061 20553 19073 20587
rect 19107 20584 19119 20587
rect 19426 20584 19432 20596
rect 19107 20556 19432 20584
rect 19107 20553 19119 20556
rect 19061 20547 19119 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20036 20556 20944 20584
rect 20036 20544 20042 20556
rect 16025 20519 16083 20525
rect 15068 20488 15424 20516
rect 15068 20476 15074 20488
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 13924 20380 13952 20408
rect 14384 20380 14412 20411
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14608 20420 14653 20448
rect 14608 20408 14614 20420
rect 14918 20408 14924 20460
rect 14976 20457 14982 20460
rect 14976 20411 14984 20457
rect 14976 20408 14982 20411
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15396 20457 15424 20488
rect 16025 20485 16037 20519
rect 16071 20485 16083 20519
rect 16025 20479 16083 20485
rect 16132 20488 19288 20516
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 15160 20420 15209 20448
rect 15160 20408 15166 20420
rect 15197 20417 15209 20420
rect 15243 20417 15255 20451
rect 15197 20411 15255 20417
rect 15381 20451 15439 20457
rect 15381 20417 15393 20451
rect 15427 20417 15439 20451
rect 15381 20411 15439 20417
rect 13004 20352 13952 20380
rect 14292 20352 14412 20380
rect 15289 20383 15347 20389
rect 12872 20343 12930 20349
rect 9600 20284 11100 20312
rect 7745 20247 7803 20253
rect 7745 20213 7757 20247
rect 7791 20213 7803 20247
rect 7745 20207 7803 20213
rect 7834 20204 7840 20256
rect 7892 20244 7898 20256
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 7892 20216 8217 20244
rect 7892 20204 7898 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 8404 20244 8432 20272
rect 9600 20244 9628 20284
rect 12342 20272 12348 20324
rect 12400 20312 12406 20324
rect 12713 20315 12771 20321
rect 12713 20312 12725 20315
rect 12400 20284 12725 20312
rect 12400 20272 12406 20284
rect 12713 20281 12725 20284
rect 12759 20281 12771 20315
rect 12713 20275 12771 20281
rect 8404 20216 9628 20244
rect 9677 20247 9735 20253
rect 8205 20207 8263 20213
rect 9677 20213 9689 20247
rect 9723 20244 9735 20247
rect 11514 20244 11520 20256
rect 9723 20216 11520 20244
rect 9723 20213 9735 20216
rect 9677 20207 9735 20213
rect 11514 20204 11520 20216
rect 11572 20204 11578 20256
rect 11698 20204 11704 20256
rect 11756 20244 11762 20256
rect 12437 20247 12495 20253
rect 12437 20244 12449 20247
rect 11756 20216 12449 20244
rect 11756 20204 11762 20216
rect 12437 20213 12449 20216
rect 12483 20213 12495 20247
rect 14292 20244 14320 20352
rect 15289 20349 15301 20383
rect 15335 20380 15347 20383
rect 16132 20380 16160 20488
rect 16206 20408 16212 20460
rect 16264 20408 16270 20460
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16301 20411 16359 20417
rect 16316 20380 16344 20411
rect 16666 20408 16672 20460
rect 16724 20408 16730 20460
rect 16850 20408 16856 20460
rect 16908 20408 16914 20460
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 17184 20420 17233 20448
rect 17184 20408 17190 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 17865 20451 17923 20457
rect 17865 20448 17877 20451
rect 17221 20411 17279 20417
rect 17328 20420 17877 20448
rect 15335 20352 16160 20380
rect 16224 20352 16344 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 14366 20272 14372 20324
rect 14424 20312 14430 20324
rect 16224 20312 16252 20352
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 16448 20352 16957 20380
rect 16448 20340 16454 20352
rect 16945 20349 16957 20352
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 17034 20340 17040 20392
rect 17092 20340 17098 20392
rect 14424 20284 16252 20312
rect 16485 20315 16543 20321
rect 14424 20272 14430 20284
rect 16485 20281 16497 20315
rect 16531 20312 16543 20315
rect 17328 20312 17356 20420
rect 17865 20417 17877 20420
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 18046 20408 18052 20460
rect 18104 20408 18110 20460
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20448 18291 20451
rect 18322 20448 18328 20460
rect 18279 20420 18328 20448
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 18690 20448 18696 20460
rect 18463 20420 18696 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19260 20457 19288 20488
rect 19352 20488 19932 20516
rect 19352 20460 19380 20488
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19334 20408 19340 20460
rect 19392 20408 19398 20460
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19904 20457 19932 20488
rect 19889 20451 19947 20457
rect 19576 20420 19621 20448
rect 19576 20408 19582 20420
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20417 20039 20451
rect 19981 20411 20039 20417
rect 18138 20340 18144 20392
rect 18196 20340 18202 20392
rect 19429 20383 19487 20389
rect 19429 20380 19441 20383
rect 18524 20352 19441 20380
rect 16531 20284 17356 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 18524 20312 18552 20352
rect 19429 20349 19441 20352
rect 19475 20380 19487 20383
rect 19996 20380 20024 20411
rect 20162 20408 20168 20460
rect 20220 20408 20226 20460
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20622 20448 20628 20460
rect 20303 20420 20628 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20916 20457 20944 20556
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21453 20587 21511 20593
rect 21453 20584 21465 20587
rect 21232 20556 21465 20584
rect 21232 20544 21238 20556
rect 21453 20553 21465 20556
rect 21499 20553 21511 20587
rect 21453 20547 21511 20553
rect 22462 20544 22468 20596
rect 22520 20584 22526 20596
rect 22557 20587 22615 20593
rect 22557 20584 22569 20587
rect 22520 20556 22569 20584
rect 22520 20544 22526 20556
rect 22557 20553 22569 20556
rect 22603 20553 22615 20587
rect 22557 20547 22615 20553
rect 24486 20544 24492 20596
rect 24544 20544 24550 20596
rect 26145 20587 26203 20593
rect 26145 20553 26157 20587
rect 26191 20584 26203 20587
rect 26326 20584 26332 20596
rect 26191 20556 26332 20584
rect 26191 20553 26203 20556
rect 26145 20547 26203 20553
rect 26326 20544 26332 20556
rect 26384 20544 26390 20596
rect 23017 20519 23075 20525
rect 23017 20516 23029 20519
rect 21008 20488 23029 20516
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20417 20959 20451
rect 20901 20411 20959 20417
rect 21008 20380 21036 20488
rect 23017 20485 23029 20488
rect 23063 20485 23075 20519
rect 24673 20519 24731 20525
rect 24673 20516 24685 20519
rect 24242 20488 24685 20516
rect 23017 20479 23075 20485
rect 24673 20485 24685 20488
rect 24719 20485 24731 20519
rect 28994 20516 29000 20528
rect 24673 20479 24731 20485
rect 26068 20488 29000 20516
rect 21082 20408 21088 20460
rect 21140 20408 21146 20460
rect 21174 20408 21180 20460
rect 21232 20408 21238 20460
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 22465 20451 22523 20457
rect 22465 20417 22477 20451
rect 22511 20448 22523 20451
rect 22554 20448 22560 20460
rect 22511 20420 22560 20448
rect 22511 20417 22523 20420
rect 22465 20411 22523 20417
rect 22554 20408 22560 20420
rect 22612 20408 22618 20460
rect 26068 20457 26096 20488
rect 28994 20476 29000 20488
rect 29052 20476 29058 20528
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20448 24823 20451
rect 26053 20451 26111 20457
rect 26053 20448 26065 20451
rect 24811 20420 26065 20448
rect 24811 20417 24823 20420
rect 24765 20411 24823 20417
rect 26053 20417 26065 20420
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 21818 20380 21824 20392
rect 19475 20352 20024 20380
rect 20824 20352 21036 20380
rect 21376 20352 21824 20380
rect 19475 20349 19487 20352
rect 19429 20343 19487 20349
rect 17552 20284 18552 20312
rect 18601 20315 18659 20321
rect 17552 20272 17558 20284
rect 18601 20281 18613 20315
rect 18647 20312 18659 20315
rect 19334 20312 19340 20324
rect 18647 20284 19340 20312
rect 18647 20281 18659 20284
rect 18601 20275 18659 20281
rect 19334 20272 19340 20284
rect 19392 20272 19398 20324
rect 19518 20272 19524 20324
rect 19576 20312 19582 20324
rect 20824 20312 20852 20352
rect 19576 20284 20852 20312
rect 19576 20272 19582 20284
rect 16206 20244 16212 20256
rect 14292 20216 16212 20244
rect 12437 20207 12495 20213
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 16301 20247 16359 20253
rect 16301 20213 16313 20247
rect 16347 20244 16359 20247
rect 16942 20244 16948 20256
rect 16347 20216 16948 20244
rect 16347 20213 16359 20216
rect 16301 20207 16359 20213
rect 16942 20204 16948 20216
rect 17000 20204 17006 20256
rect 17405 20247 17463 20253
rect 17405 20213 17417 20247
rect 17451 20244 17463 20247
rect 17862 20244 17868 20256
rect 17451 20216 17868 20244
rect 17451 20213 17463 20216
rect 17405 20207 17463 20213
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 19705 20247 19763 20253
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 19794 20244 19800 20256
rect 19751 20216 19800 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 21376 20244 21404 20352
rect 21818 20340 21824 20352
rect 21876 20380 21882 20392
rect 21876 20352 22094 20380
rect 21876 20340 21882 20352
rect 20772 20216 21404 20244
rect 22066 20244 22094 20352
rect 22186 20340 22192 20392
rect 22244 20380 22250 20392
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 22244 20352 22753 20380
rect 22244 20340 22250 20352
rect 22741 20349 22753 20352
rect 22787 20349 22799 20383
rect 24780 20380 24808 20411
rect 27522 20408 27528 20460
rect 27580 20408 27586 20460
rect 24946 20380 24952 20392
rect 22741 20343 22799 20349
rect 22848 20352 24952 20380
rect 22554 20272 22560 20324
rect 22612 20312 22618 20324
rect 22848 20312 22876 20352
rect 24946 20340 24952 20352
rect 25004 20340 25010 20392
rect 27617 20383 27675 20389
rect 27617 20349 27629 20383
rect 27663 20380 27675 20383
rect 27706 20380 27712 20392
rect 27663 20352 27712 20380
rect 27663 20349 27675 20352
rect 27617 20343 27675 20349
rect 27706 20340 27712 20352
rect 27764 20340 27770 20392
rect 29086 20312 29092 20324
rect 22612 20284 22876 20312
rect 24044 20284 29092 20312
rect 22612 20272 22618 20284
rect 24044 20244 24072 20284
rect 29086 20272 29092 20284
rect 29144 20272 29150 20324
rect 22066 20216 24072 20244
rect 27801 20247 27859 20253
rect 20772 20204 20778 20216
rect 27801 20213 27813 20247
rect 27847 20244 27859 20247
rect 27890 20244 27896 20256
rect 27847 20216 27896 20244
rect 27847 20213 27859 20216
rect 27801 20207 27859 20213
rect 27890 20204 27896 20216
rect 27948 20204 27954 20256
rect 1104 20154 29716 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 29716 20154
rect 1104 20080 29716 20102
rect 4525 20043 4583 20049
rect 4525 20009 4537 20043
rect 4571 20040 4583 20043
rect 4798 20040 4804 20052
rect 4571 20012 4804 20040
rect 4571 20009 4583 20012
rect 4525 20003 4583 20009
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 6178 20000 6184 20052
rect 6236 20000 6242 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 7984 20012 8432 20040
rect 7984 20000 7990 20012
rect 4890 19972 4896 19984
rect 2792 19944 4896 19972
rect 2792 19913 2820 19944
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 5905 19975 5963 19981
rect 5905 19941 5917 19975
rect 5951 19972 5963 19975
rect 6454 19972 6460 19984
rect 5951 19944 6460 19972
rect 5951 19941 5963 19944
rect 5905 19935 5963 19941
rect 6454 19932 6460 19944
rect 6512 19932 6518 19984
rect 6730 19932 6736 19984
rect 6788 19972 6794 19984
rect 8404 19972 8432 20012
rect 8938 20000 8944 20052
rect 8996 20040 9002 20052
rect 9033 20043 9091 20049
rect 9033 20040 9045 20043
rect 8996 20012 9045 20040
rect 8996 20000 9002 20012
rect 9033 20009 9045 20012
rect 9079 20040 9091 20043
rect 9858 20040 9864 20052
rect 9079 20012 9864 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 11238 20040 11244 20052
rect 9968 20012 11244 20040
rect 9968 19972 9996 20012
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 16666 20040 16672 20052
rect 11572 20012 11928 20040
rect 11572 20000 11578 20012
rect 6788 19944 8340 19972
rect 8404 19944 9996 19972
rect 10045 19975 10103 19981
rect 6788 19932 6794 19944
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19873 2835 19907
rect 2777 19867 2835 19873
rect 6638 19864 6644 19916
rect 6696 19864 6702 19916
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 900 19808 1501 19836
rect 900 19796 906 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1489 19799 1547 19805
rect 1670 19796 1676 19848
rect 1728 19796 1734 19848
rect 2866 19796 2872 19848
rect 2924 19836 2930 19848
rect 4062 19836 4068 19848
rect 2924 19808 4068 19836
rect 2924 19796 2930 19808
rect 4062 19796 4068 19808
rect 4120 19836 4126 19848
rect 4433 19839 4491 19845
rect 4433 19836 4445 19839
rect 4120 19808 4445 19836
rect 4120 19796 4126 19808
rect 4433 19805 4445 19808
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 5810 19796 5816 19848
rect 5868 19796 5874 19848
rect 6270 19796 6276 19848
rect 6328 19796 6334 19848
rect 6362 19796 6368 19848
rect 6420 19796 6426 19848
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6748 19845 6776 19932
rect 7466 19864 7472 19916
rect 7524 19864 7530 19916
rect 7834 19904 7840 19916
rect 7668 19876 7840 19904
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19805 6791 19839
rect 6733 19799 6791 19805
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19836 6975 19839
rect 7282 19836 7288 19848
rect 6963 19808 7288 19836
rect 6963 19805 6975 19808
rect 6917 19799 6975 19805
rect 2685 19771 2743 19777
rect 2685 19737 2697 19771
rect 2731 19768 2743 19771
rect 3418 19768 3424 19780
rect 2731 19740 3424 19768
rect 2731 19737 2743 19740
rect 2685 19731 2743 19737
rect 3418 19728 3424 19740
rect 3476 19768 3482 19780
rect 5828 19768 5856 19796
rect 3476 19740 5856 19768
rect 3476 19728 3482 19740
rect 6454 19728 6460 19780
rect 6512 19768 6518 19780
rect 6748 19768 6776 19799
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7668 19845 7696 19876
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7653 19839 7711 19845
rect 7653 19805 7665 19839
rect 7699 19805 7711 19839
rect 7653 19799 7711 19805
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8110 19836 8116 19848
rect 7791 19808 8116 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 6512 19740 6776 19768
rect 7392 19768 7420 19799
rect 8110 19796 8116 19808
rect 8168 19796 8174 19848
rect 8202 19796 8208 19848
rect 8260 19796 8266 19848
rect 8312 19836 8340 19944
rect 10045 19941 10057 19975
rect 10091 19972 10103 19975
rect 11330 19972 11336 19984
rect 10091 19944 11336 19972
rect 10091 19941 10103 19944
rect 10045 19935 10103 19941
rect 11330 19932 11336 19944
rect 11388 19972 11394 19984
rect 11388 19944 11652 19972
rect 11388 19932 11394 19944
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 8536 19876 8984 19904
rect 8536 19864 8542 19876
rect 8956 19845 8984 19876
rect 9490 19864 9496 19916
rect 9548 19904 9554 19916
rect 11624 19913 11652 19944
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 9548 19876 10272 19904
rect 9548 19864 9554 19876
rect 8389 19839 8447 19845
rect 8389 19836 8401 19839
rect 8312 19808 8401 19836
rect 8389 19805 8401 19808
rect 8435 19805 8447 19839
rect 8389 19799 8447 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 8573 19799 8631 19805
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 7392 19740 8248 19768
rect 6512 19728 6518 19740
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2225 19703 2283 19709
rect 2225 19700 2237 19703
rect 1728 19672 2237 19700
rect 1728 19660 1734 19672
rect 2225 19669 2237 19672
rect 2271 19669 2283 19703
rect 2225 19663 2283 19669
rect 2590 19660 2596 19712
rect 2648 19660 2654 19712
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 7064 19672 7113 19700
rect 7064 19660 7070 19672
rect 7101 19669 7113 19672
rect 7147 19669 7159 19703
rect 7101 19663 7159 19669
rect 7926 19660 7932 19712
rect 7984 19660 7990 19712
rect 8018 19660 8024 19712
rect 8076 19660 8082 19712
rect 8220 19700 8248 19740
rect 8294 19728 8300 19780
rect 8352 19728 8358 19780
rect 8588 19768 8616 19799
rect 9766 19796 9772 19848
rect 9824 19836 9830 19848
rect 9953 19839 10011 19845
rect 9953 19836 9965 19839
rect 9824 19808 9965 19836
rect 9824 19796 9830 19808
rect 9953 19805 9965 19808
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10244 19845 10272 19876
rect 10980 19876 11437 19904
rect 10137 19839 10195 19845
rect 10137 19836 10149 19839
rect 10100 19808 10149 19836
rect 10100 19796 10106 19808
rect 10137 19805 10149 19808
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 10413 19839 10471 19845
rect 10413 19805 10425 19839
rect 10459 19805 10471 19839
rect 10413 19799 10471 19805
rect 9122 19768 9128 19780
rect 8588 19740 9128 19768
rect 9122 19728 9128 19740
rect 9180 19768 9186 19780
rect 9490 19768 9496 19780
rect 9180 19740 9496 19768
rect 9180 19728 9186 19740
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 9674 19728 9680 19780
rect 9732 19768 9738 19780
rect 10428 19768 10456 19799
rect 10686 19796 10692 19848
rect 10744 19796 10750 19848
rect 10778 19796 10784 19848
rect 10836 19796 10842 19848
rect 10980 19845 11008 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 11698 19864 11704 19916
rect 11756 19864 11762 19916
rect 11900 19913 11928 20012
rect 14752 20012 16672 20040
rect 14752 19984 14780 20012
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 16758 20000 16764 20052
rect 16816 20040 16822 20052
rect 16853 20043 16911 20049
rect 16853 20040 16865 20043
rect 16816 20012 16865 20040
rect 16816 20000 16822 20012
rect 16853 20009 16865 20012
rect 16899 20009 16911 20043
rect 16853 20003 16911 20009
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 17310 20040 17316 20052
rect 17000 20012 17316 20040
rect 17000 20000 17006 20012
rect 17310 20000 17316 20012
rect 17368 20000 17374 20052
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 18196 20012 18337 20040
rect 18196 20000 18202 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 18325 20003 18383 20009
rect 19426 20000 19432 20052
rect 19484 20040 19490 20052
rect 19886 20040 19892 20052
rect 19484 20012 19892 20040
rect 19484 20000 19490 20012
rect 19886 20000 19892 20012
rect 19944 20040 19950 20052
rect 20625 20043 20683 20049
rect 19944 20012 20576 20040
rect 19944 20000 19950 20012
rect 14734 19972 14740 19984
rect 14568 19944 14740 19972
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 9732 19740 10456 19768
rect 9732 19728 9738 19740
rect 10594 19728 10600 19780
rect 10652 19768 10658 19780
rect 11057 19771 11115 19777
rect 11057 19768 11069 19771
rect 10652 19740 11069 19768
rect 10652 19728 10658 19740
rect 11057 19737 11069 19740
rect 11103 19737 11115 19771
rect 11057 19731 11115 19737
rect 11164 19768 11192 19799
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11296 19808 11805 19836
rect 11296 19796 11302 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 11793 19799 11851 19805
rect 12406 19808 12725 19836
rect 11974 19768 11980 19780
rect 11164 19740 11980 19768
rect 8754 19700 8760 19712
rect 8220 19672 8760 19700
rect 8754 19660 8760 19672
rect 8812 19660 8818 19712
rect 10413 19703 10471 19709
rect 10413 19669 10425 19703
rect 10459 19700 10471 19703
rect 11164 19700 11192 19740
rect 11974 19728 11980 19740
rect 12032 19728 12038 19780
rect 10459 19672 11192 19700
rect 11333 19703 11391 19709
rect 10459 19669 10471 19672
rect 10413 19663 10471 19669
rect 11333 19669 11345 19703
rect 11379 19700 11391 19703
rect 12406 19700 12434 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13354 19836 13360 19848
rect 13035 19808 13360 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 14568 19845 14596 19944
rect 14734 19932 14740 19944
rect 14792 19932 14798 19984
rect 15289 19975 15347 19981
rect 15289 19941 15301 19975
rect 15335 19941 15347 19975
rect 15289 19935 15347 19941
rect 15304 19904 15332 19935
rect 16206 19932 16212 19984
rect 16264 19972 16270 19984
rect 17126 19972 17132 19984
rect 16264 19944 17132 19972
rect 16264 19932 16270 19944
rect 17126 19932 17132 19944
rect 17184 19932 17190 19984
rect 18046 19932 18052 19984
rect 18104 19972 18110 19984
rect 18417 19975 18475 19981
rect 18417 19972 18429 19975
rect 18104 19944 18429 19972
rect 18104 19932 18110 19944
rect 18417 19941 18429 19944
rect 18463 19941 18475 19975
rect 19705 19975 19763 19981
rect 19705 19972 19717 19975
rect 18417 19935 18475 19941
rect 18800 19944 19717 19972
rect 18800 19904 18828 19944
rect 19705 19941 19717 19944
rect 19751 19941 19763 19975
rect 19705 19935 19763 19941
rect 19794 19932 19800 19984
rect 19852 19932 19858 19984
rect 14660 19876 14872 19904
rect 15304 19876 18828 19904
rect 14660 19845 14688 19876
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19805 14703 19839
rect 14645 19799 14703 19805
rect 14738 19839 14796 19845
rect 14738 19805 14750 19839
rect 14784 19805 14796 19839
rect 14738 19799 14796 19805
rect 14752 19768 14780 19799
rect 14568 19740 14780 19768
rect 14568 19712 14596 19740
rect 11379 19672 12434 19700
rect 12805 19703 12863 19709
rect 11379 19669 11391 19672
rect 11333 19663 11391 19669
rect 12805 19669 12817 19703
rect 12851 19700 12863 19703
rect 12986 19700 12992 19712
rect 12851 19672 12992 19700
rect 12851 19669 12863 19672
rect 12805 19663 12863 19669
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 13170 19660 13176 19712
rect 13228 19660 13234 19712
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 14550 19700 14556 19712
rect 14507 19672 14556 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 14844 19700 14872 19876
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20548 19904 20576 20012
rect 20625 20009 20637 20043
rect 20671 20040 20683 20043
rect 21726 20040 21732 20052
rect 20671 20012 21732 20040
rect 20671 20009 20683 20012
rect 20625 20003 20683 20009
rect 21726 20000 21732 20012
rect 21784 20000 21790 20052
rect 26697 20043 26755 20049
rect 26697 20009 26709 20043
rect 26743 20040 26755 20043
rect 26743 20012 27292 20040
rect 26743 20009 26755 20012
rect 26697 20003 26755 20009
rect 21174 19932 21180 19984
rect 21232 19972 21238 19984
rect 21910 19972 21916 19984
rect 21232 19944 21916 19972
rect 21232 19932 21238 19944
rect 21910 19932 21916 19944
rect 21968 19932 21974 19984
rect 21545 19907 21603 19913
rect 20548 19876 21220 19904
rect 14918 19796 14924 19848
rect 14976 19796 14982 19848
rect 15102 19796 15108 19848
rect 15160 19845 15166 19848
rect 15160 19836 15168 19845
rect 15160 19808 15205 19836
rect 15160 19799 15168 19808
rect 15160 19796 15166 19799
rect 15562 19796 15568 19848
rect 15620 19796 15626 19848
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17402 19836 17408 19848
rect 16991 19808 17408 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17402 19796 17408 19808
rect 17460 19836 17466 19848
rect 17586 19836 17592 19848
rect 17460 19808 17592 19836
rect 17460 19796 17466 19808
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 17681 19839 17739 19845
rect 17681 19805 17693 19839
rect 17727 19805 17739 19839
rect 17681 19799 17739 19805
rect 15010 19728 15016 19780
rect 15068 19768 15074 19780
rect 15473 19771 15531 19777
rect 15473 19768 15485 19771
rect 15068 19740 15485 19768
rect 15068 19728 15074 19740
rect 15473 19737 15485 19740
rect 15519 19737 15531 19771
rect 15473 19731 15531 19737
rect 16666 19728 16672 19780
rect 16724 19768 16730 19780
rect 17494 19768 17500 19780
rect 16724 19740 17500 19768
rect 16724 19728 16730 19740
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 17696 19768 17724 19799
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 18138 19796 18144 19848
rect 18196 19796 18202 19848
rect 18322 19796 18328 19848
rect 18380 19836 18386 19848
rect 18601 19839 18659 19845
rect 18601 19836 18613 19839
rect 18380 19808 18613 19836
rect 18380 19796 18386 19808
rect 18601 19805 18613 19808
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 18748 19808 18936 19836
rect 18748 19796 18754 19808
rect 17954 19768 17960 19780
rect 17696 19740 17960 19768
rect 17954 19728 17960 19740
rect 18012 19768 18018 19780
rect 18230 19768 18236 19780
rect 18012 19740 18236 19768
rect 18012 19728 18018 19740
rect 18230 19728 18236 19740
rect 18288 19728 18294 19780
rect 18782 19728 18788 19780
rect 18840 19728 18846 19780
rect 18908 19768 18936 19808
rect 18966 19796 18972 19848
rect 19024 19796 19030 19848
rect 19610 19796 19616 19848
rect 19668 19845 19674 19848
rect 19668 19839 19683 19845
rect 19671 19805 19683 19839
rect 19668 19799 19683 19805
rect 19668 19796 19674 19799
rect 19886 19796 19892 19848
rect 19944 19796 19950 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 19242 19768 19248 19780
rect 18908 19740 19248 19768
rect 19242 19728 19248 19740
rect 19300 19728 19306 19780
rect 19429 19771 19487 19777
rect 19429 19737 19441 19771
rect 19475 19768 19487 19771
rect 20364 19768 20392 19799
rect 20438 19796 20444 19848
rect 20496 19796 20502 19848
rect 21082 19796 21088 19848
rect 21140 19796 21146 19848
rect 21192 19845 21220 19876
rect 21545 19873 21557 19907
rect 21591 19904 21603 19907
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 21591 19876 22109 19904
rect 21591 19873 21603 19876
rect 21545 19867 21603 19873
rect 22097 19873 22109 19876
rect 22143 19904 22155 19907
rect 22278 19904 22284 19916
rect 22143 19876 22284 19904
rect 22143 19873 22155 19876
rect 22097 19867 22155 19873
rect 22278 19864 22284 19876
rect 22336 19864 22342 19916
rect 23290 19864 23296 19916
rect 23348 19904 23354 19916
rect 24949 19907 25007 19913
rect 24949 19904 24961 19907
rect 23348 19876 24961 19904
rect 23348 19864 23354 19876
rect 24949 19873 24961 19876
rect 24995 19904 25007 19907
rect 26234 19904 26240 19916
rect 24995 19876 26240 19904
rect 24995 19873 25007 19876
rect 24949 19867 25007 19873
rect 26234 19864 26240 19876
rect 26292 19864 26298 19916
rect 26878 19864 26884 19916
rect 26936 19904 26942 19916
rect 27264 19913 27292 20012
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 29365 20043 29423 20049
rect 29365 20040 29377 20043
rect 27580 20012 29377 20040
rect 27580 20000 27586 20012
rect 29365 20009 29377 20012
rect 29411 20009 29423 20043
rect 29365 20003 29423 20009
rect 27157 19907 27215 19913
rect 27157 19904 27169 19907
rect 26936 19876 27169 19904
rect 26936 19864 26942 19876
rect 27157 19873 27169 19876
rect 27203 19873 27215 19907
rect 27157 19867 27215 19873
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19904 27307 19907
rect 27338 19904 27344 19916
rect 27295 19876 27344 19904
rect 27295 19873 27307 19876
rect 27249 19867 27307 19873
rect 27338 19864 27344 19876
rect 27396 19864 27402 19916
rect 21177 19839 21235 19845
rect 21177 19805 21189 19839
rect 21223 19805 21235 19839
rect 21177 19799 21235 19805
rect 21358 19796 21364 19848
rect 21416 19836 21422 19848
rect 21821 19839 21879 19845
rect 21821 19836 21833 19839
rect 21416 19808 21833 19836
rect 21416 19796 21422 19808
rect 21821 19805 21833 19808
rect 21867 19805 21879 19839
rect 21821 19799 21879 19805
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22189 19839 22247 19845
rect 22189 19836 22201 19839
rect 22066 19808 22201 19836
rect 19475 19740 20392 19768
rect 21453 19771 21511 19777
rect 19475 19737 19487 19740
rect 19429 19731 19487 19737
rect 21453 19737 21465 19771
rect 21499 19768 21511 19771
rect 22066 19768 22094 19808
rect 22189 19805 22201 19808
rect 22235 19836 22247 19839
rect 22830 19836 22836 19848
rect 22235 19808 22836 19836
rect 22235 19805 22247 19808
rect 22189 19799 22247 19805
rect 22830 19796 22836 19808
rect 22888 19796 22894 19848
rect 26970 19796 26976 19848
rect 27028 19796 27034 19848
rect 27065 19839 27123 19845
rect 27065 19805 27077 19839
rect 27111 19836 27123 19839
rect 27540 19836 27568 20000
rect 27614 19864 27620 19916
rect 27672 19864 27678 19916
rect 27890 19864 27896 19916
rect 27948 19864 27954 19916
rect 27111 19808 27568 19836
rect 27111 19805 27123 19808
rect 27065 19799 27123 19805
rect 27264 19780 27292 19808
rect 21499 19740 22094 19768
rect 21499 19737 21511 19740
rect 21453 19731 21511 19737
rect 21836 19712 21864 19740
rect 25130 19728 25136 19780
rect 25188 19768 25194 19780
rect 25225 19771 25283 19777
rect 25225 19768 25237 19771
rect 25188 19740 25237 19768
rect 25188 19728 25194 19740
rect 25225 19737 25237 19740
rect 25271 19737 25283 19771
rect 25225 19731 25283 19737
rect 25958 19728 25964 19780
rect 26016 19728 26022 19780
rect 27246 19728 27252 19780
rect 27304 19728 27310 19780
rect 28902 19728 28908 19780
rect 28960 19728 28966 19780
rect 20806 19700 20812 19712
rect 14844 19672 20812 19700
rect 20806 19660 20812 19672
rect 20864 19700 20870 19712
rect 20901 19703 20959 19709
rect 20901 19700 20913 19703
rect 20864 19672 20913 19700
rect 20864 19660 20870 19672
rect 20901 19669 20913 19672
rect 20947 19669 20959 19703
rect 20901 19663 20959 19669
rect 21634 19660 21640 19712
rect 21692 19660 21698 19712
rect 21818 19660 21824 19712
rect 21876 19660 21882 19712
rect 26786 19660 26792 19712
rect 26844 19660 26850 19712
rect 1104 19610 29716 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 29716 19610
rect 1104 19536 29716 19558
rect 7466 19456 7472 19508
rect 7524 19456 7530 19508
rect 8662 19456 8668 19508
rect 8720 19456 8726 19508
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 9946 19499 10004 19505
rect 9946 19465 9958 19499
rect 9992 19496 10004 19499
rect 10594 19496 10600 19508
rect 9992 19468 10600 19496
rect 9992 19465 10004 19468
rect 9946 19459 10004 19465
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 10873 19499 10931 19505
rect 10873 19496 10885 19499
rect 10744 19468 10885 19496
rect 10744 19456 10750 19468
rect 10873 19465 10885 19468
rect 10919 19465 10931 19499
rect 10873 19459 10931 19465
rect 12161 19499 12219 19505
rect 12161 19465 12173 19499
rect 12207 19496 12219 19499
rect 12989 19499 13047 19505
rect 12207 19468 12480 19496
rect 12207 19465 12219 19468
rect 12161 19459 12219 19465
rect 1670 19388 1676 19440
rect 1728 19388 1734 19440
rect 3418 19388 3424 19440
rect 3476 19388 3482 19440
rect 5169 19431 5227 19437
rect 5169 19397 5181 19431
rect 5215 19428 5227 19431
rect 5534 19428 5540 19440
rect 5215 19400 5540 19428
rect 5215 19397 5227 19400
rect 5169 19391 5227 19397
rect 5534 19388 5540 19400
rect 5592 19388 5598 19440
rect 8018 19428 8024 19440
rect 6932 19400 8024 19428
rect 6932 19372 6960 19400
rect 8018 19388 8024 19400
rect 8076 19388 8082 19440
rect 8680 19428 8708 19456
rect 9122 19428 9128 19440
rect 8496 19400 9128 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 3786 19320 3792 19372
rect 3844 19360 3850 19372
rect 3844 19332 4752 19360
rect 3844 19320 3850 19332
rect 4724 19233 4752 19332
rect 5074 19320 5080 19372
rect 5132 19320 5138 19372
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 6914 19320 6920 19372
rect 6972 19320 6978 19372
rect 7006 19320 7012 19372
rect 7064 19320 7070 19372
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19360 7343 19363
rect 7374 19360 7380 19372
rect 7331 19332 7380 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7374 19320 7380 19332
rect 7432 19360 7438 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 7432 19332 8125 19360
rect 7432 19320 7438 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8297 19363 8355 19369
rect 8297 19360 8309 19363
rect 8113 19323 8171 19329
rect 8220 19332 8309 19360
rect 4890 19252 4896 19304
rect 4948 19292 4954 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 4948 19264 5273 19292
rect 4948 19252 4954 19264
rect 5261 19261 5273 19264
rect 5307 19261 5319 19295
rect 5261 19255 5319 19261
rect 7101 19295 7159 19301
rect 7101 19261 7113 19295
rect 7147 19292 7159 19295
rect 7742 19292 7748 19304
rect 7147 19264 7748 19292
rect 7147 19261 7159 19264
rect 7101 19255 7159 19261
rect 4709 19227 4767 19233
rect 4709 19193 4721 19227
rect 4755 19193 4767 19227
rect 4709 19187 4767 19193
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 7116 19224 7144 19255
rect 7742 19252 7748 19264
rect 7800 19292 7806 19304
rect 8220 19292 8248 19332
rect 8297 19329 8309 19332
rect 8343 19329 8355 19363
rect 8297 19323 8355 19329
rect 8386 19320 8392 19372
rect 8444 19320 8450 19372
rect 8496 19369 8524 19400
rect 9122 19388 9128 19400
rect 9180 19388 9186 19440
rect 9858 19388 9864 19440
rect 9916 19388 9922 19440
rect 10612 19428 10640 19456
rect 11793 19431 11851 19437
rect 11793 19428 11805 19431
rect 10612 19400 11805 19428
rect 11793 19397 11805 19400
rect 11839 19397 11851 19431
rect 11793 19391 11851 19397
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 8941 19363 8999 19369
rect 8941 19360 8953 19363
rect 8720 19332 8953 19360
rect 8720 19320 8726 19332
rect 8941 19329 8953 19332
rect 8987 19329 8999 19363
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 8941 19323 8999 19329
rect 9232 19332 9321 19360
rect 7800 19264 8248 19292
rect 8404 19292 8432 19320
rect 9232 19301 9260 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9456 19332 9505 19360
rect 9456 19320 9462 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19329 9827 19363
rect 9769 19323 9827 19329
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 10502 19360 10508 19372
rect 10091 19332 10508 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 8404 19264 9229 19292
rect 7800 19252 7806 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9784 19292 9812 19323
rect 10502 19320 10508 19332
rect 10560 19360 10566 19372
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 10560 19332 10793 19360
rect 10560 19320 10566 19332
rect 10781 19329 10793 19332
rect 10827 19329 10839 19363
rect 10781 19323 10839 19329
rect 10962 19320 10968 19372
rect 11020 19360 11026 19372
rect 12452 19369 12480 19468
rect 12989 19465 13001 19499
rect 13035 19496 13047 19499
rect 15194 19496 15200 19508
rect 13035 19468 15200 19496
rect 13035 19465 13047 19468
rect 12989 19459 13047 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 17184 19468 17724 19496
rect 17184 19456 17190 19468
rect 12621 19431 12679 19437
rect 12621 19397 12633 19431
rect 12667 19428 12679 19431
rect 13262 19428 13268 19440
rect 12667 19400 13268 19428
rect 12667 19397 12679 19400
rect 12621 19391 12679 19397
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 14090 19388 14096 19440
rect 14148 19428 14154 19440
rect 17310 19428 17316 19440
rect 14148 19400 14504 19428
rect 14148 19388 14154 19400
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11020 19332 11897 19360
rect 11020 19320 11026 19332
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 12002 19363 12060 19369
rect 12002 19329 12014 19363
rect 12048 19360 12060 19363
rect 12437 19363 12495 19369
rect 12048 19332 12296 19360
rect 12048 19329 12060 19332
rect 12002 19323 12060 19329
rect 9858 19292 9864 19304
rect 9784 19264 9864 19292
rect 9217 19255 9275 19261
rect 9858 19252 9864 19264
rect 9916 19292 9922 19304
rect 10226 19292 10232 19304
rect 9916 19264 10232 19292
rect 9916 19252 9922 19264
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 11514 19252 11520 19304
rect 11572 19252 11578 19304
rect 12268 19292 12296 19332
rect 12437 19329 12449 19363
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12713 19363 12771 19369
rect 12713 19329 12725 19363
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 12805 19363 12863 19369
rect 12805 19329 12817 19363
rect 12851 19360 12863 19363
rect 13170 19360 13176 19372
rect 12851 19332 13176 19360
rect 12851 19329 12863 19332
rect 12805 19323 12863 19329
rect 12342 19292 12348 19304
rect 12268 19264 12348 19292
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 7064 19196 7144 19224
rect 9401 19227 9459 19233
rect 7064 19184 7070 19196
rect 9401 19193 9413 19227
rect 9447 19224 9459 19227
rect 12158 19224 12164 19236
rect 9447 19196 12164 19224
rect 9447 19193 9459 19196
rect 9401 19187 9459 19193
rect 12158 19184 12164 19196
rect 12216 19224 12222 19236
rect 12728 19224 12756 19323
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14476 19369 14504 19400
rect 16868 19400 17316 19428
rect 16868 19372 16896 19400
rect 17310 19388 17316 19400
rect 17368 19388 17374 19440
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 14240 19332 14289 19360
rect 14240 19320 14246 19332
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 14734 19360 14740 19372
rect 14507 19332 14740 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 14829 19363 14887 19369
rect 14829 19329 14841 19363
rect 14875 19360 14887 19363
rect 15010 19360 15016 19372
rect 14875 19332 15016 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 15010 19320 15016 19332
rect 15068 19320 15074 19372
rect 16850 19320 16856 19372
rect 16908 19320 16914 19372
rect 16942 19320 16948 19372
rect 17000 19320 17006 19372
rect 17221 19363 17279 19369
rect 17221 19329 17233 19363
rect 17267 19360 17279 19363
rect 17494 19360 17500 19372
rect 17267 19332 17500 19360
rect 17267 19329 17279 19332
rect 17221 19323 17279 19329
rect 17494 19320 17500 19332
rect 17552 19320 17558 19372
rect 17696 19369 17724 19468
rect 18230 19456 18236 19508
rect 18288 19456 18294 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20438 19496 20444 19508
rect 19843 19468 20444 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20438 19456 20444 19468
rect 20496 19456 20502 19508
rect 20622 19456 20628 19508
rect 20680 19456 20686 19508
rect 20815 19499 20873 19505
rect 20815 19496 20827 19499
rect 20732 19468 20827 19496
rect 17862 19388 17868 19440
rect 17920 19388 17926 19440
rect 17954 19388 17960 19440
rect 18012 19428 18018 19440
rect 18874 19428 18880 19440
rect 18012 19400 18880 19428
rect 18012 19388 18018 19400
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 19426 19388 19432 19440
rect 19484 19388 19490 19440
rect 19886 19388 19892 19440
rect 19944 19428 19950 19440
rect 20732 19428 20760 19468
rect 20815 19465 20827 19468
rect 20861 19465 20873 19499
rect 20815 19459 20873 19465
rect 20901 19499 20959 19505
rect 20901 19465 20913 19499
rect 20947 19496 20959 19499
rect 21634 19496 21640 19508
rect 20947 19468 21640 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 22830 19456 22836 19508
rect 22888 19496 22894 19508
rect 24673 19499 24731 19505
rect 24673 19496 24685 19499
rect 22888 19468 24685 19496
rect 22888 19456 22894 19468
rect 24673 19465 24685 19468
rect 24719 19465 24731 19499
rect 24673 19459 24731 19465
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 25958 19456 25964 19508
rect 26016 19456 26022 19508
rect 27246 19456 27252 19508
rect 27304 19456 27310 19508
rect 27338 19456 27344 19508
rect 27396 19456 27402 19508
rect 27706 19456 27712 19508
rect 27764 19456 27770 19508
rect 28902 19456 28908 19508
rect 28960 19456 28966 19508
rect 19944 19400 20760 19428
rect 19944 19388 19950 19400
rect 21358 19388 21364 19440
rect 21416 19388 21422 19440
rect 23290 19428 23296 19440
rect 22940 19400 23296 19428
rect 17681 19363 17739 19369
rect 17681 19329 17693 19363
rect 17727 19329 17739 19363
rect 17681 19323 17739 19329
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19360 18107 19363
rect 18322 19360 18328 19372
rect 18095 19332 18328 19360
rect 18095 19329 18107 19332
rect 18049 19323 18107 19329
rect 18322 19320 18328 19332
rect 18380 19320 18386 19372
rect 18966 19320 18972 19372
rect 19024 19360 19030 19372
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 19024 19332 19257 19360
rect 19024 19320 19030 19332
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 14550 19252 14556 19304
rect 14608 19252 14614 19304
rect 14642 19252 14648 19304
rect 14700 19252 14706 19304
rect 16758 19252 16764 19304
rect 16816 19292 16822 19304
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16816 19264 17141 19292
rect 16816 19252 16822 19264
rect 17129 19261 17141 19264
rect 17175 19261 17187 19295
rect 19260 19292 19288 19323
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19392 19332 19533 19360
rect 19392 19320 19398 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 19702 19320 19708 19372
rect 19760 19360 19766 19372
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19760 19332 19993 19360
rect 19760 19320 19766 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 19981 19323 20039 19329
rect 20070 19320 20076 19372
rect 20128 19360 20134 19372
rect 20257 19363 20315 19369
rect 20128 19332 20173 19360
rect 20128 19320 20134 19332
rect 20257 19329 20269 19363
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 19260 19264 20208 19292
rect 17129 19255 17187 19261
rect 12216 19196 12756 19224
rect 12216 19184 12222 19196
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 16022 19224 16028 19236
rect 14332 19196 16028 19224
rect 14332 19184 14338 19196
rect 16022 19184 16028 19196
rect 16080 19224 16086 19236
rect 16942 19224 16948 19236
rect 16080 19196 16948 19224
rect 16080 19184 16086 19196
rect 16942 19184 16948 19196
rect 17000 19184 17006 19236
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 9122 19116 9128 19168
rect 9180 19116 9186 19168
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15286 19156 15292 19168
rect 15059 19128 15292 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 15896 19128 16681 19156
rect 15896 19116 15902 19128
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 20180 19156 20208 19264
rect 20272 19224 20300 19323
rect 20346 19320 20352 19372
rect 20404 19320 20410 19372
rect 20487 19363 20545 19369
rect 20487 19329 20499 19363
rect 20533 19360 20545 19363
rect 20622 19360 20628 19372
rect 20533 19332 20628 19360
rect 20533 19329 20545 19332
rect 20487 19323 20545 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 20717 19363 20775 19369
rect 20717 19329 20729 19363
rect 20763 19360 20775 19363
rect 20806 19360 20812 19372
rect 20763 19332 20812 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 20990 19320 20996 19372
rect 21048 19320 21054 19372
rect 21450 19360 21456 19372
rect 21192 19332 21456 19360
rect 21192 19224 21220 19332
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 22940 19369 22968 19400
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 24857 19431 24915 19437
rect 24857 19428 24869 19431
rect 24426 19400 24869 19428
rect 24857 19397 24869 19400
rect 24903 19397 24915 19431
rect 24857 19391 24915 19397
rect 29270 19388 29276 19440
rect 29328 19388 29334 19440
rect 22925 19363 22983 19369
rect 22925 19329 22937 19363
rect 22971 19329 22983 19363
rect 22925 19323 22983 19329
rect 24670 19320 24676 19372
rect 24728 19360 24734 19372
rect 24946 19360 24952 19372
rect 24728 19332 24952 19360
rect 24728 19320 24734 19332
rect 24946 19320 24952 19332
rect 25004 19360 25010 19372
rect 25869 19363 25927 19369
rect 25869 19360 25881 19363
rect 25004 19332 25881 19360
rect 25004 19320 25010 19332
rect 25869 19329 25881 19332
rect 25915 19360 25927 19363
rect 26234 19360 26240 19372
rect 25915 19332 26240 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 27154 19320 27160 19372
rect 27212 19360 27218 19372
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 27212 19332 27629 19360
rect 27212 19320 27218 19332
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 27801 19363 27859 19369
rect 27801 19329 27813 19363
rect 27847 19329 27859 19363
rect 27801 19323 27859 19329
rect 22462 19252 22468 19304
rect 22520 19292 22526 19304
rect 23201 19295 23259 19301
rect 23201 19292 23213 19295
rect 22520 19264 23213 19292
rect 22520 19252 22526 19264
rect 23201 19261 23213 19264
rect 23247 19261 23259 19295
rect 23201 19255 23259 19261
rect 25593 19295 25651 19301
rect 25593 19261 25605 19295
rect 25639 19292 25651 19295
rect 26050 19292 26056 19304
rect 25639 19264 26056 19292
rect 25639 19261 25651 19264
rect 25593 19255 25651 19261
rect 26050 19252 26056 19264
rect 26108 19292 26114 19304
rect 26973 19295 27031 19301
rect 26973 19292 26985 19295
rect 26108 19264 26985 19292
rect 26108 19252 26114 19264
rect 26973 19261 26985 19264
rect 27019 19261 27031 19295
rect 27816 19292 27844 19323
rect 28994 19320 29000 19372
rect 29052 19320 29058 19372
rect 26973 19255 27031 19261
rect 27540 19264 27844 19292
rect 27540 19236 27568 19264
rect 20272 19196 21220 19224
rect 25317 19227 25375 19233
rect 25317 19193 25329 19227
rect 25363 19224 25375 19227
rect 26786 19224 26792 19236
rect 25363 19196 26792 19224
rect 25363 19193 25375 19196
rect 25317 19187 25375 19193
rect 26786 19184 26792 19196
rect 26844 19184 26850 19236
rect 26878 19184 26884 19236
rect 26936 19224 26942 19236
rect 27522 19224 27528 19236
rect 26936 19196 27528 19224
rect 26936 19184 26942 19196
rect 27522 19184 27528 19196
rect 27580 19184 27586 19236
rect 21082 19156 21088 19168
rect 20180 19128 21088 19156
rect 16669 19119 16727 19125
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 29181 19159 29239 19165
rect 29181 19125 29193 19159
rect 29227 19156 29239 19159
rect 29638 19156 29644 19168
rect 29227 19128 29644 19156
rect 29227 19125 29239 19128
rect 29181 19119 29239 19125
rect 29638 19116 29644 19128
rect 29696 19116 29702 19168
rect 1104 19066 29716 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 29716 19066
rect 1104 18992 29716 19014
rect 2409 18955 2467 18961
rect 2409 18921 2421 18955
rect 2455 18952 2467 18955
rect 2774 18952 2780 18964
rect 2455 18924 2780 18952
rect 2455 18921 2467 18924
rect 2409 18915 2467 18921
rect 2774 18912 2780 18924
rect 2832 18912 2838 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3200 18924 3801 18952
rect 3200 18912 3206 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 4890 18952 4896 18964
rect 4396 18924 4896 18952
rect 4396 18912 4402 18924
rect 4890 18912 4896 18924
rect 4948 18912 4954 18964
rect 6454 18952 6460 18964
rect 5000 18924 6460 18952
rect 5000 18884 5028 18924
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 6825 18955 6883 18961
rect 6825 18921 6837 18955
rect 6871 18952 6883 18955
rect 6914 18952 6920 18964
rect 6871 18924 6920 18952
rect 6871 18921 6883 18924
rect 6825 18915 6883 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 7190 18912 7196 18964
rect 7248 18912 7254 18964
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 7340 18924 7389 18952
rect 7340 18912 7346 18924
rect 7377 18921 7389 18924
rect 7423 18952 7435 18955
rect 9490 18952 9496 18964
rect 7423 18924 9496 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 10502 18912 10508 18964
rect 10560 18912 10566 18964
rect 16850 18952 16856 18964
rect 14200 18924 16856 18952
rect 2746 18856 5028 18884
rect 1673 18819 1731 18825
rect 1673 18785 1685 18819
rect 1719 18816 1731 18819
rect 2746 18816 2774 18856
rect 5074 18844 5080 18896
rect 5132 18844 5138 18896
rect 5718 18884 5724 18896
rect 5460 18856 5724 18884
rect 1719 18788 2774 18816
rect 3973 18819 4031 18825
rect 1719 18785 1731 18788
rect 1673 18779 1731 18785
rect 3973 18785 3985 18819
rect 4019 18816 4031 18819
rect 4154 18816 4160 18828
rect 4019 18788 4160 18816
rect 4019 18785 4031 18788
rect 3973 18779 4031 18785
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 5460 18825 5488 18856
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 8662 18884 8668 18896
rect 7024 18856 8668 18884
rect 4617 18819 4675 18825
rect 4617 18816 4629 18819
rect 4304 18788 4629 18816
rect 4304 18776 4310 18788
rect 4617 18785 4629 18788
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18785 5227 18819
rect 5169 18779 5227 18785
rect 5445 18819 5503 18825
rect 5445 18785 5457 18819
rect 5491 18785 5503 18819
rect 5445 18779 5503 18785
rect 842 18708 848 18760
rect 900 18748 906 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 900 18720 1409 18748
rect 900 18708 906 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18748 2375 18751
rect 2866 18748 2872 18760
rect 2363 18720 2872 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 4062 18708 4068 18760
rect 4120 18708 4126 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18748 4862 18760
rect 5184 18748 5212 18779
rect 5626 18776 5632 18828
rect 5684 18816 5690 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 5684 18788 6837 18816
rect 5684 18776 5690 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 4856 18720 5212 18748
rect 4856 18708 4862 18720
rect 5534 18708 5540 18760
rect 5592 18708 5598 18760
rect 7024 18757 7052 18856
rect 8662 18844 8668 18856
rect 8720 18844 8726 18896
rect 9585 18887 9643 18893
rect 9585 18853 9597 18887
rect 9631 18884 9643 18887
rect 9674 18884 9680 18896
rect 9631 18856 9680 18884
rect 9631 18853 9643 18856
rect 9585 18847 9643 18853
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 10045 18887 10103 18893
rect 10045 18853 10057 18887
rect 10091 18884 10103 18887
rect 10962 18884 10968 18896
rect 10091 18856 10968 18884
rect 10091 18853 10103 18856
rect 10045 18847 10103 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 14200 18884 14228 18924
rect 16850 18912 16856 18924
rect 16908 18912 16914 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18509 18955 18567 18961
rect 18509 18952 18521 18955
rect 18196 18924 18521 18952
rect 18196 18912 18202 18924
rect 18509 18921 18521 18924
rect 18555 18921 18567 18955
rect 18509 18915 18567 18921
rect 18601 18955 18659 18961
rect 18601 18921 18613 18955
rect 18647 18952 18659 18955
rect 18690 18952 18696 18964
rect 18647 18924 18696 18952
rect 18647 18921 18659 18924
rect 18601 18915 18659 18921
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 21082 18912 21088 18964
rect 21140 18952 21146 18964
rect 21269 18955 21327 18961
rect 21269 18952 21281 18955
rect 21140 18924 21281 18952
rect 21140 18912 21146 18924
rect 21269 18921 21281 18924
rect 21315 18921 21327 18955
rect 21269 18915 21327 18921
rect 22462 18912 22468 18964
rect 22520 18912 22526 18964
rect 14108 18856 14228 18884
rect 8202 18816 8208 18828
rect 8036 18788 8208 18816
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 7098 18708 7104 18760
rect 7156 18748 7162 18760
rect 7282 18748 7288 18760
rect 7156 18720 7288 18748
rect 7156 18708 7162 18720
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 8036 18757 8064 18788
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18785 8355 18819
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8297 18779 8355 18785
rect 8404 18788 9045 18816
rect 8021 18751 8079 18757
rect 8021 18748 8033 18751
rect 7524 18720 8033 18748
rect 7524 18708 7530 18720
rect 8021 18717 8033 18720
rect 8067 18717 8079 18751
rect 8021 18711 8079 18717
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18717 8171 18751
rect 8113 18711 8171 18717
rect 3878 18640 3884 18692
rect 3936 18680 3942 18692
rect 4338 18680 4344 18692
rect 3936 18652 4344 18680
rect 3936 18640 3942 18652
rect 4338 18640 4344 18652
rect 4396 18640 4402 18692
rect 4430 18640 4436 18692
rect 4488 18680 4494 18692
rect 4614 18680 4620 18692
rect 4488 18652 4620 18680
rect 4488 18640 4494 18652
rect 4614 18640 4620 18652
rect 4672 18680 4678 18692
rect 6270 18680 6276 18692
rect 4672 18652 6276 18680
rect 4672 18640 4678 18652
rect 6270 18640 6276 18652
rect 6328 18640 6334 18692
rect 6549 18683 6607 18689
rect 6549 18649 6561 18683
rect 6595 18680 6607 18683
rect 6730 18680 6736 18692
rect 6595 18652 6736 18680
rect 6595 18649 6607 18652
rect 6549 18643 6607 18649
rect 6730 18640 6736 18652
rect 6788 18680 6794 18692
rect 7837 18683 7895 18689
rect 7837 18680 7849 18683
rect 6788 18652 7849 18680
rect 6788 18640 6794 18652
rect 7837 18649 7849 18652
rect 7883 18649 7895 18683
rect 7837 18643 7895 18649
rect 8128 18612 8156 18711
rect 8312 18680 8340 18779
rect 8404 18760 8432 18788
rect 9033 18785 9045 18788
rect 9079 18785 9091 18819
rect 10137 18819 10195 18825
rect 10137 18816 10149 18819
rect 9033 18779 9091 18785
rect 9692 18788 10149 18816
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 8938 18708 8944 18760
rect 8996 18708 9002 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9692 18748 9720 18788
rect 10137 18785 10149 18788
rect 10183 18785 10195 18819
rect 10137 18779 10195 18785
rect 9548 18720 9720 18748
rect 9548 18708 9554 18720
rect 9766 18708 9772 18760
rect 9824 18708 9830 18760
rect 9858 18708 9864 18760
rect 9916 18708 9922 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 9122 18680 9128 18692
rect 8312 18652 9128 18680
rect 9122 18640 9128 18652
rect 9180 18640 9186 18692
rect 9674 18640 9680 18692
rect 9732 18680 9738 18692
rect 10134 18680 10140 18692
rect 9732 18652 10140 18680
rect 9732 18640 9738 18652
rect 10134 18640 10140 18652
rect 10192 18680 10198 18692
rect 10336 18680 10364 18711
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 14108 18757 14136 18856
rect 14366 18844 14372 18896
rect 14424 18884 14430 18896
rect 15289 18887 15347 18893
rect 14424 18856 15148 18884
rect 14424 18844 14430 18856
rect 14182 18776 14188 18828
rect 14240 18816 14246 18828
rect 14240 18788 15056 18816
rect 14240 18776 14246 18788
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 10468 18720 14105 18748
rect 10468 18708 10474 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 14366 18708 14372 18760
rect 14424 18708 14430 18760
rect 14461 18751 14519 18757
rect 14461 18717 14473 18751
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 10192 18652 10364 18680
rect 14476 18680 14504 18711
rect 14550 18708 14556 18760
rect 14608 18748 14614 18760
rect 14645 18751 14703 18757
rect 14645 18748 14657 18751
rect 14608 18720 14657 18748
rect 14608 18708 14614 18720
rect 14645 18717 14657 18720
rect 14691 18717 14703 18751
rect 14645 18711 14703 18717
rect 14734 18708 14740 18760
rect 14792 18708 14798 18760
rect 15028 18757 15056 18788
rect 15120 18757 15148 18856
rect 15289 18853 15301 18887
rect 15335 18853 15347 18887
rect 15289 18847 15347 18853
rect 15013 18751 15071 18757
rect 15013 18717 15025 18751
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 15105 18751 15163 18757
rect 15105 18717 15117 18751
rect 15151 18717 15163 18751
rect 15304 18748 15332 18847
rect 17126 18844 17132 18896
rect 17184 18884 17190 18896
rect 18874 18884 18880 18896
rect 17184 18856 18276 18884
rect 17184 18844 17190 18856
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 17770 18816 17776 18828
rect 17267 18788 17776 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 17770 18776 17776 18788
rect 17828 18816 17834 18828
rect 17828 18788 18092 18816
rect 17828 18776 17834 18788
rect 15657 18751 15715 18757
rect 15657 18748 15669 18751
rect 15304 18720 15669 18748
rect 15105 18711 15163 18717
rect 15657 18717 15669 18720
rect 15703 18717 15715 18751
rect 15657 18711 15715 18717
rect 15838 18708 15844 18760
rect 15896 18708 15902 18760
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17126 18748 17132 18760
rect 17083 18720 17132 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 17402 18708 17408 18760
rect 17460 18708 17466 18760
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17552 18720 17601 18748
rect 17552 18708 17558 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17589 18711 17647 18717
rect 17678 18708 17684 18760
rect 17736 18748 17742 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17736 18720 17877 18748
rect 17736 18708 17742 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 17954 18708 17960 18760
rect 18012 18708 18018 18760
rect 18064 18757 18092 18788
rect 18248 18757 18276 18856
rect 18524 18856 18880 18884
rect 18524 18825 18552 18856
rect 18874 18844 18880 18856
rect 18932 18884 18938 18896
rect 20346 18884 20352 18896
rect 18932 18856 20352 18884
rect 18932 18844 18938 18856
rect 20346 18844 20352 18856
rect 20404 18884 20410 18896
rect 20404 18856 22232 18884
rect 20404 18844 20410 18856
rect 18509 18819 18567 18825
rect 18509 18785 18521 18819
rect 18555 18785 18567 18819
rect 20070 18816 20076 18828
rect 18509 18779 18567 18785
rect 18616 18788 20076 18816
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18616 18748 18644 18788
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 21634 18776 21640 18828
rect 21692 18816 21698 18828
rect 22097 18819 22155 18825
rect 22097 18816 22109 18819
rect 21692 18788 22109 18816
rect 21692 18776 21698 18788
rect 22097 18785 22109 18788
rect 22143 18785 22155 18819
rect 22097 18779 22155 18785
rect 22204 18760 22232 18856
rect 27709 18819 27767 18825
rect 27709 18785 27721 18819
rect 27755 18816 27767 18819
rect 27755 18788 28028 18816
rect 27755 18785 27767 18788
rect 27709 18779 27767 18785
rect 18279 18720 18644 18748
rect 18693 18751 18751 18757
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18693 18717 18705 18751
rect 18739 18748 18751 18751
rect 18966 18748 18972 18760
rect 18739 18720 18972 18748
rect 18739 18717 18751 18720
rect 18693 18711 18751 18717
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19978 18748 19984 18760
rect 19392 18720 19984 18748
rect 19392 18708 19398 18720
rect 19978 18708 19984 18720
rect 20036 18748 20042 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 20036 18720 20361 18748
rect 20036 18708 20042 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 20349 18711 20407 18717
rect 21358 18708 21364 18760
rect 21416 18708 21422 18760
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 22741 18751 22799 18757
rect 22741 18748 22753 18751
rect 22244 18720 22753 18748
rect 22244 18708 22250 18720
rect 22741 18717 22753 18720
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 22830 18708 22836 18760
rect 22888 18708 22894 18760
rect 27798 18708 27804 18760
rect 27856 18708 27862 18760
rect 28000 18757 28028 18788
rect 29086 18776 29092 18828
rect 29144 18776 29150 18828
rect 27985 18751 28043 18757
rect 27985 18717 27997 18751
rect 28031 18717 28043 18751
rect 27985 18711 28043 18717
rect 29362 18708 29368 18760
rect 29420 18708 29426 18760
rect 14476 18652 15240 18680
rect 10192 18640 10198 18652
rect 8294 18612 8300 18624
rect 8128 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 10318 18612 10324 18624
rect 8352 18584 10324 18612
rect 8352 18572 8358 18584
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 14918 18572 14924 18624
rect 14976 18572 14982 18624
rect 15212 18612 15240 18652
rect 15286 18640 15292 18692
rect 15344 18640 15350 18692
rect 17328 18680 17356 18708
rect 15764 18652 17080 18680
rect 17328 18652 17908 18680
rect 15764 18612 15792 18652
rect 17052 18624 17080 18652
rect 15212 18584 15792 18612
rect 15841 18615 15899 18621
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 16758 18612 16764 18624
rect 15887 18584 16764 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 16850 18572 16856 18624
rect 16908 18572 16914 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 17092 18584 17693 18612
rect 17092 18572 17098 18584
rect 17681 18581 17693 18584
rect 17727 18581 17739 18615
rect 17880 18612 17908 18652
rect 18322 18640 18328 18692
rect 18380 18680 18386 18692
rect 18874 18680 18880 18692
rect 18380 18652 18880 18680
rect 18380 18640 18386 18652
rect 18874 18640 18880 18652
rect 18932 18640 18938 18692
rect 26786 18640 26792 18692
rect 26844 18680 26850 18692
rect 27154 18680 27160 18692
rect 26844 18652 27160 18680
rect 26844 18640 26850 18652
rect 27154 18640 27160 18652
rect 27212 18680 27218 18692
rect 27341 18683 27399 18689
rect 27341 18680 27353 18683
rect 27212 18652 27353 18680
rect 27212 18640 27218 18652
rect 27341 18649 27353 18652
rect 27387 18649 27399 18683
rect 27341 18643 27399 18649
rect 27522 18640 27528 18692
rect 27580 18640 27586 18692
rect 20257 18615 20315 18621
rect 20257 18612 20269 18615
rect 17880 18584 20269 18612
rect 17681 18575 17739 18581
rect 20257 18581 20269 18584
rect 20303 18581 20315 18615
rect 20257 18575 20315 18581
rect 27890 18572 27896 18624
rect 27948 18612 27954 18624
rect 28169 18615 28227 18621
rect 28169 18612 28181 18615
rect 27948 18584 28181 18612
rect 27948 18572 27954 18584
rect 28169 18581 28181 18584
rect 28215 18581 28227 18615
rect 28169 18575 28227 18581
rect 1104 18522 29716 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 29716 18522
rect 1104 18448 29716 18470
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2590 18408 2596 18420
rect 2547 18380 2596 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 4065 18411 4123 18417
rect 4065 18377 4077 18411
rect 4111 18408 4123 18411
rect 4430 18408 4436 18420
rect 4111 18380 4436 18408
rect 4111 18377 4123 18380
rect 4065 18371 4123 18377
rect 4430 18368 4436 18380
rect 4488 18368 4494 18420
rect 11054 18408 11060 18420
rect 10796 18380 11060 18408
rect 1673 18343 1731 18349
rect 1673 18309 1685 18343
rect 1719 18340 1731 18343
rect 10410 18340 10416 18352
rect 1719 18312 10416 18340
rect 1719 18309 1731 18312
rect 1673 18303 1731 18309
rect 10410 18300 10416 18312
rect 10468 18300 10474 18352
rect 10796 18349 10824 18380
rect 11054 18368 11060 18380
rect 11112 18408 11118 18420
rect 12066 18408 12072 18420
rect 11112 18380 12072 18408
rect 11112 18368 11118 18380
rect 12066 18368 12072 18380
rect 12124 18408 12130 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 12124 18380 13553 18408
rect 12124 18368 12130 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 13541 18371 13599 18377
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15381 18411 15439 18417
rect 15381 18408 15393 18411
rect 15344 18380 15393 18408
rect 15344 18368 15350 18380
rect 15381 18377 15393 18380
rect 15427 18377 15439 18411
rect 15381 18371 15439 18377
rect 17494 18368 17500 18420
rect 17552 18368 17558 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 18598 18408 18604 18420
rect 18380 18380 18604 18408
rect 18380 18368 18386 18380
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 20070 18368 20076 18420
rect 20128 18408 20134 18420
rect 20990 18408 20996 18420
rect 20128 18380 20996 18408
rect 20128 18368 20134 18380
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 21416 18380 25053 18408
rect 21416 18368 21422 18380
rect 15194 18349 15200 18352
rect 10781 18343 10839 18349
rect 10781 18309 10793 18343
rect 10827 18309 10839 18343
rect 13817 18343 13875 18349
rect 13817 18340 13829 18343
rect 13294 18312 13829 18340
rect 10781 18303 10839 18309
rect 13817 18309 13829 18312
rect 13863 18309 13875 18343
rect 13817 18303 13875 18309
rect 15172 18343 15200 18349
rect 15172 18309 15184 18343
rect 15172 18303 15200 18309
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 1854 18272 1860 18284
rect 1811 18244 1860 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 1854 18232 1860 18244
rect 1912 18232 1918 18284
rect 2130 18232 2136 18284
rect 2188 18232 2194 18284
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 3973 18275 4031 18281
rect 3973 18272 3985 18275
rect 3200 18244 3985 18272
rect 3200 18232 3206 18244
rect 3973 18241 3985 18244
rect 4019 18241 4031 18275
rect 3973 18235 4031 18241
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 3326 18204 3332 18216
rect 2271 18176 3332 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 3988 18204 4016 18235
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 4212 18244 4261 18272
rect 4212 18232 4218 18244
rect 4249 18241 4261 18244
rect 4295 18272 4307 18275
rect 4614 18272 4620 18284
rect 4295 18244 4620 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 5258 18232 5264 18284
rect 5316 18272 5322 18284
rect 5442 18272 5448 18284
rect 5316 18244 5448 18272
rect 5316 18232 5322 18244
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18272 10287 18275
rect 10796 18272 10824 18303
rect 15194 18300 15200 18303
rect 15252 18300 15258 18352
rect 16850 18340 16856 18352
rect 15304 18312 16856 18340
rect 10275 18244 10824 18272
rect 10275 18241 10287 18244
rect 10229 18235 10287 18241
rect 10962 18232 10968 18284
rect 11020 18232 11026 18284
rect 11790 18232 11796 18284
rect 11848 18232 11854 18284
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14274 18272 14280 18284
rect 13955 18244 14280 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 5718 18204 5724 18216
rect 3988 18176 5724 18204
rect 5718 18164 5724 18176
rect 5776 18164 5782 18216
rect 10318 18164 10324 18216
rect 10376 18204 10382 18216
rect 10870 18204 10876 18216
rect 10376 18176 10876 18204
rect 10376 18164 10382 18176
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 12066 18164 12072 18216
rect 12124 18164 12130 18216
rect 15304 18213 15332 18312
rect 16850 18300 16856 18312
rect 16908 18340 16914 18352
rect 16945 18343 17003 18349
rect 16945 18340 16957 18343
rect 16908 18312 16957 18340
rect 16908 18300 16914 18312
rect 16945 18309 16957 18312
rect 16991 18309 17003 18343
rect 16945 18303 17003 18309
rect 15488 18244 15792 18272
rect 15289 18207 15347 18213
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15289 18167 15347 18173
rect 4246 18096 4252 18148
rect 4304 18096 4310 18148
rect 5350 18096 5356 18148
rect 5408 18136 5414 18148
rect 5534 18136 5540 18148
rect 5408 18108 5540 18136
rect 5408 18096 5414 18108
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 8938 18096 8944 18148
rect 8996 18136 9002 18148
rect 8996 18108 10824 18136
rect 8996 18096 9002 18108
rect 10796 18080 10824 18108
rect 14918 18096 14924 18148
rect 14976 18136 14982 18148
rect 15488 18136 15516 18244
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18173 15715 18207
rect 15764 18204 15792 18244
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 15896 18244 16313 18272
rect 15896 18232 15902 18244
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 15764 18176 16037 18204
rect 15657 18167 15715 18173
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 16025 18167 16083 18173
rect 16684 18204 16712 18235
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 16816 18244 16861 18272
rect 16816 18232 16822 18244
rect 17034 18232 17040 18284
rect 17092 18232 17098 18284
rect 17175 18275 17233 18281
rect 17175 18241 17187 18275
rect 17221 18272 17233 18275
rect 17512 18272 17540 18368
rect 18064 18312 18736 18340
rect 17221 18244 17540 18272
rect 17221 18241 17233 18244
rect 17175 18235 17233 18241
rect 17678 18232 17684 18284
rect 17736 18232 17742 18284
rect 17773 18275 17831 18281
rect 17773 18241 17785 18275
rect 17819 18272 17831 18275
rect 17954 18272 17960 18284
rect 17819 18244 17960 18272
rect 17819 18241 17831 18244
rect 17773 18235 17831 18241
rect 17954 18232 17960 18244
rect 18012 18232 18018 18284
rect 18064 18281 18092 18312
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 18322 18232 18328 18284
rect 18380 18232 18386 18284
rect 18414 18232 18420 18284
rect 18472 18232 18478 18284
rect 18708 18281 18736 18312
rect 18509 18275 18567 18281
rect 18509 18241 18521 18275
rect 18555 18272 18567 18275
rect 18693 18275 18751 18281
rect 18555 18244 18644 18272
rect 18555 18241 18567 18244
rect 18509 18235 18567 18241
rect 16684 18176 18184 18204
rect 14976 18108 15516 18136
rect 15672 18136 15700 18167
rect 15749 18139 15807 18145
rect 15749 18136 15761 18139
rect 15672 18108 15761 18136
rect 14976 18096 14982 18108
rect 15749 18105 15761 18108
rect 15795 18105 15807 18139
rect 15749 18099 15807 18105
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10468 18040 10609 18068
rect 10468 18028 10474 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 10778 18028 10784 18080
rect 10836 18068 10842 18080
rect 12618 18068 12624 18080
rect 10836 18040 12624 18068
rect 10836 18028 10842 18040
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15654 18068 15660 18080
rect 15059 18040 15660 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15654 18028 15660 18040
rect 15712 18028 15718 18080
rect 16209 18071 16267 18077
rect 16209 18037 16221 18071
rect 16255 18068 16267 18071
rect 16684 18068 16712 18176
rect 16850 18096 16856 18148
rect 16908 18136 16914 18148
rect 17678 18136 17684 18148
rect 16908 18108 17684 18136
rect 16908 18096 16914 18108
rect 17678 18096 17684 18108
rect 17736 18096 17742 18148
rect 18156 18145 18184 18176
rect 18141 18139 18199 18145
rect 18141 18105 18153 18139
rect 18187 18105 18199 18139
rect 18141 18099 18199 18105
rect 16255 18040 16712 18068
rect 16255 18037 16267 18040
rect 16209 18031 16267 18037
rect 17310 18028 17316 18080
rect 17368 18028 17374 18080
rect 17957 18071 18015 18077
rect 17957 18037 17969 18071
rect 18003 18068 18015 18071
rect 18506 18068 18512 18080
rect 18003 18040 18512 18068
rect 18003 18037 18015 18040
rect 17957 18031 18015 18037
rect 18506 18028 18512 18040
rect 18564 18068 18570 18080
rect 18616 18068 18644 18244
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 18966 18272 18972 18284
rect 18739 18244 18972 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 21174 18272 21180 18284
rect 21131 18244 21180 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 21266 18232 21272 18284
rect 21324 18272 21330 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 21324 18244 21373 18272
rect 21324 18232 21330 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18241 21511 18275
rect 21453 18235 21511 18241
rect 21468 18204 21496 18235
rect 21542 18232 21548 18284
rect 21600 18272 21606 18284
rect 21637 18275 21695 18281
rect 21637 18272 21649 18275
rect 21600 18244 21649 18272
rect 21600 18232 21606 18244
rect 21637 18241 21649 18244
rect 21683 18272 21695 18275
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21683 18244 21833 18272
rect 21683 18241 21695 18244
rect 21637 18235 21695 18241
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 21910 18232 21916 18284
rect 21968 18232 21974 18284
rect 22848 18281 22876 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 27522 18368 27528 18420
rect 27580 18408 27586 18420
rect 29365 18411 29423 18417
rect 29365 18408 29377 18411
rect 27580 18380 29377 18408
rect 27580 18368 27586 18380
rect 29365 18377 29377 18380
rect 29411 18377 29423 18411
rect 29365 18371 29423 18377
rect 24578 18300 24584 18352
rect 24636 18300 24642 18352
rect 27890 18300 27896 18352
rect 27948 18300 27954 18352
rect 28902 18300 28908 18352
rect 28960 18300 28966 18352
rect 22097 18275 22155 18281
rect 22097 18241 22109 18275
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 22189 18275 22247 18281
rect 22189 18241 22201 18275
rect 22235 18272 22247 18275
rect 22833 18275 22891 18281
rect 22235 18244 22324 18272
rect 22235 18241 22247 18244
rect 22189 18235 22247 18241
rect 21468 18176 22048 18204
rect 21634 18096 21640 18148
rect 21692 18096 21698 18148
rect 22020 18080 22048 18176
rect 22112 18136 22140 18235
rect 22186 18136 22192 18148
rect 22112 18108 22192 18136
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 18782 18068 18788 18080
rect 18564 18040 18788 18068
rect 18564 18028 18570 18040
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 22002 18028 22008 18080
rect 22060 18068 22066 18080
rect 22296 18068 22324 18244
rect 22833 18241 22845 18275
rect 22879 18241 22891 18275
rect 22833 18235 22891 18241
rect 23290 18232 23296 18284
rect 23348 18232 23354 18284
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 22373 18207 22431 18213
rect 22373 18173 22385 18207
rect 22419 18204 22431 18207
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22419 18176 22753 18204
rect 22419 18173 22431 18176
rect 22373 18167 22431 18173
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 23569 18207 23627 18213
rect 23569 18204 23581 18207
rect 22741 18167 22799 18173
rect 23216 18176 23581 18204
rect 23216 18145 23244 18176
rect 23569 18173 23581 18176
rect 23615 18173 23627 18207
rect 23569 18167 23627 18173
rect 25038 18164 25044 18216
rect 25096 18204 25102 18216
rect 25225 18207 25283 18213
rect 25225 18204 25237 18207
rect 25096 18176 25237 18204
rect 25096 18164 25102 18176
rect 25225 18173 25237 18176
rect 25271 18173 25283 18207
rect 25332 18204 25360 18235
rect 26234 18232 26240 18284
rect 26292 18232 26298 18284
rect 27614 18232 27620 18284
rect 27672 18232 27678 18284
rect 26326 18204 26332 18216
rect 25332 18176 26332 18204
rect 25225 18167 25283 18173
rect 26326 18164 26332 18176
rect 26384 18164 26390 18216
rect 23201 18139 23259 18145
rect 23201 18105 23213 18139
rect 23247 18105 23259 18139
rect 23201 18099 23259 18105
rect 22060 18040 22324 18068
rect 22060 18028 22066 18040
rect 25498 18028 25504 18080
rect 25556 18068 25562 18080
rect 25593 18071 25651 18077
rect 25593 18068 25605 18071
rect 25556 18040 25605 18068
rect 25556 18028 25562 18040
rect 25593 18037 25605 18040
rect 25639 18037 25651 18071
rect 25593 18031 25651 18037
rect 26234 18028 26240 18080
rect 26292 18068 26298 18080
rect 26329 18071 26387 18077
rect 26329 18068 26341 18071
rect 26292 18040 26341 18068
rect 26292 18028 26298 18040
rect 26329 18037 26341 18040
rect 26375 18037 26387 18071
rect 26329 18031 26387 18037
rect 1104 17978 29716 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 29716 17978
rect 1104 17904 29716 17926
rect 2130 17824 2136 17876
rect 2188 17864 2194 17876
rect 2317 17867 2375 17873
rect 2317 17864 2329 17867
rect 2188 17836 2329 17864
rect 2188 17824 2194 17836
rect 2317 17833 2329 17836
rect 2363 17833 2375 17867
rect 2317 17827 2375 17833
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 3418 17864 3424 17876
rect 2556 17836 3424 17864
rect 2556 17824 2562 17836
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 3789 17867 3847 17873
rect 3789 17833 3801 17867
rect 3835 17864 3847 17867
rect 4062 17864 4068 17876
rect 3835 17836 4068 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 6270 17864 6276 17876
rect 5828 17836 6276 17864
rect 2593 17799 2651 17805
rect 2593 17765 2605 17799
rect 2639 17796 2651 17799
rect 4154 17796 4160 17808
rect 2639 17768 4160 17796
rect 2639 17765 2651 17768
rect 2593 17759 2651 17765
rect 2608 17728 2636 17759
rect 4154 17756 4160 17768
rect 4212 17796 4218 17808
rect 5169 17799 5227 17805
rect 4212 17768 5053 17796
rect 4212 17756 4218 17768
rect 2240 17700 2636 17728
rect 3421 17731 3479 17737
rect 2240 17669 2268 17700
rect 3421 17697 3433 17731
rect 3467 17728 3479 17731
rect 3973 17731 4031 17737
rect 3973 17728 3985 17731
rect 3467 17700 3985 17728
rect 3467 17697 3479 17700
rect 3421 17691 3479 17697
rect 3973 17697 3985 17700
rect 4019 17697 4031 17731
rect 3973 17691 4031 17697
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4338 17728 4344 17740
rect 4111 17700 4344 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4338 17688 4344 17700
rect 4396 17728 4402 17740
rect 4396 17700 4568 17728
rect 4396 17688 4402 17700
rect 2225 17663 2283 17669
rect 2225 17629 2237 17663
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 2424 17592 2452 17623
rect 2498 17620 2504 17672
rect 2556 17620 2562 17672
rect 2700 17669 2820 17670
rect 2678 17663 2820 17669
rect 2678 17629 2690 17663
rect 2724 17660 2820 17663
rect 2961 17663 3019 17669
rect 2724 17642 2912 17660
rect 2724 17629 2736 17642
rect 2792 17632 2912 17642
rect 2678 17623 2736 17629
rect 2777 17595 2835 17601
rect 2777 17592 2789 17595
rect 2424 17564 2789 17592
rect 2777 17561 2789 17564
rect 2823 17561 2835 17595
rect 2884 17592 2912 17632
rect 2961 17629 2973 17663
rect 3007 17660 3019 17663
rect 3007 17632 3280 17660
rect 3007 17629 3019 17632
rect 2961 17623 3019 17629
rect 3142 17592 3148 17604
rect 2884 17564 3148 17592
rect 2777 17555 2835 17561
rect 2792 17524 2820 17555
rect 3142 17552 3148 17564
rect 3200 17552 3206 17604
rect 3252 17592 3280 17632
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17629 3571 17663
rect 3513 17623 3571 17629
rect 3418 17592 3424 17604
rect 3252 17564 3424 17592
rect 3418 17552 3424 17564
rect 3476 17552 3482 17604
rect 3528 17592 3556 17623
rect 3786 17620 3792 17672
rect 3844 17660 3850 17672
rect 4154 17660 4160 17672
rect 3844 17632 4160 17660
rect 3844 17620 3850 17632
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 4246 17620 4252 17672
rect 4304 17620 4310 17672
rect 4540 17669 4568 17700
rect 4798 17688 4804 17740
rect 4856 17688 4862 17740
rect 5025 17737 5053 17768
rect 5169 17765 5181 17799
rect 5215 17796 5227 17799
rect 5350 17796 5356 17808
rect 5215 17768 5356 17796
rect 5215 17765 5227 17768
rect 5169 17759 5227 17765
rect 5350 17756 5356 17768
rect 5408 17756 5414 17808
rect 5010 17731 5068 17737
rect 5010 17697 5022 17731
rect 5056 17697 5068 17731
rect 5010 17691 5068 17697
rect 5718 17688 5724 17740
rect 5776 17688 5782 17740
rect 4525 17663 4583 17669
rect 4525 17629 4537 17663
rect 4571 17660 4583 17663
rect 5629 17663 5687 17669
rect 4571 17632 5304 17660
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 4893 17595 4951 17601
rect 4893 17592 4905 17595
rect 3528 17564 4905 17592
rect 3528 17524 3556 17564
rect 4893 17561 4905 17564
rect 4939 17561 4951 17595
rect 4893 17555 4951 17561
rect 2792 17496 3556 17524
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 4246 17524 4252 17536
rect 3936 17496 4252 17524
rect 3936 17484 3942 17496
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 5276 17533 5304 17632
rect 5629 17629 5641 17663
rect 5675 17660 5687 17663
rect 5828 17660 5856 17836
rect 6270 17824 6276 17836
rect 6328 17864 6334 17876
rect 8113 17867 8171 17873
rect 8113 17864 8125 17867
rect 6328 17836 8125 17864
rect 6328 17824 6334 17836
rect 8113 17833 8125 17836
rect 8159 17833 8171 17867
rect 8294 17864 8300 17876
rect 8113 17827 8171 17833
rect 8220 17836 8300 17864
rect 8220 17796 8248 17836
rect 8294 17824 8300 17836
rect 8352 17864 8358 17876
rect 8938 17864 8944 17876
rect 8352 17836 8944 17864
rect 8352 17824 8358 17836
rect 8938 17824 8944 17836
rect 8996 17824 9002 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 10744 17836 10793 17864
rect 10744 17824 10750 17836
rect 10781 17833 10793 17836
rect 10827 17864 10839 17867
rect 11793 17867 11851 17873
rect 10827 17836 11376 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 8036 17768 8248 17796
rect 8573 17799 8631 17805
rect 8036 17737 8064 17768
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 11348 17796 11376 17836
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 12066 17864 12072 17876
rect 11839 17836 12072 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 16577 17867 16635 17873
rect 16577 17833 16589 17867
rect 16623 17864 16635 17867
rect 18322 17864 18328 17876
rect 16623 17836 18328 17864
rect 16623 17833 16635 17836
rect 16577 17827 16635 17833
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 22097 17867 22155 17873
rect 22097 17864 22109 17867
rect 21968 17836 22109 17864
rect 21968 17824 21974 17836
rect 22097 17833 22109 17836
rect 22143 17833 22155 17867
rect 22097 17827 22155 17833
rect 24489 17867 24547 17873
rect 24489 17833 24501 17867
rect 24535 17864 24547 17867
rect 24578 17864 24584 17876
rect 24535 17836 24584 17864
rect 24535 17833 24547 17836
rect 24489 17827 24547 17833
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 28813 17867 28871 17873
rect 28813 17833 28825 17867
rect 28859 17864 28871 17867
rect 28902 17864 28908 17876
rect 28859 17836 28908 17864
rect 28859 17833 28871 17836
rect 28813 17827 28871 17833
rect 28902 17824 28908 17836
rect 28960 17824 28966 17876
rect 12526 17796 12532 17808
rect 8619 17768 11284 17796
rect 11348 17768 12532 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17697 8079 17731
rect 8021 17691 8079 17697
rect 5675 17632 5856 17660
rect 5675 17629 5687 17632
rect 5629 17623 5687 17629
rect 5994 17620 6000 17672
rect 6052 17620 6058 17672
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7616 17632 8309 17660
rect 7616 17620 7622 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17660 8447 17663
rect 8478 17660 8484 17672
rect 8435 17632 8484 17660
rect 8435 17629 8447 17632
rect 8389 17623 8447 17629
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8956 17669 8984 17768
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17728 10747 17731
rect 11054 17728 11060 17740
rect 10735 17700 11060 17728
rect 10735 17697 10747 17700
rect 10689 17691 10747 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9171 17632 10732 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 6273 17595 6331 17601
rect 6273 17561 6285 17595
rect 6319 17561 6331 17595
rect 6273 17555 6331 17561
rect 5261 17527 5319 17533
rect 5261 17493 5273 17527
rect 5307 17493 5319 17527
rect 6288 17524 6316 17555
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 7834 17552 7840 17604
rect 7892 17592 7898 17604
rect 8113 17595 8171 17601
rect 8113 17592 8125 17595
rect 7892 17564 8125 17592
rect 7892 17552 7898 17564
rect 8113 17561 8125 17564
rect 8159 17561 8171 17595
rect 9140 17592 9168 17623
rect 8113 17555 8171 17561
rect 8496 17564 9168 17592
rect 7098 17524 7104 17536
rect 6288 17496 7104 17524
rect 5261 17487 5319 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 8496 17524 8524 17564
rect 9858 17552 9864 17604
rect 9916 17592 9922 17604
rect 10505 17595 10563 17601
rect 10505 17592 10517 17595
rect 9916 17564 10517 17592
rect 9916 17552 9922 17564
rect 10505 17561 10517 17564
rect 10551 17561 10563 17595
rect 10704 17592 10732 17632
rect 10778 17620 10784 17672
rect 10836 17620 10842 17672
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11256 17669 11284 17768
rect 12526 17756 12532 17768
rect 12584 17796 12590 17808
rect 13722 17796 13728 17808
rect 12584 17768 13728 17796
rect 12584 17756 12590 17768
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 17954 17756 17960 17808
rect 18012 17796 18018 17808
rect 18690 17796 18696 17808
rect 18012 17768 18696 17796
rect 18012 17756 18018 17768
rect 18690 17756 18696 17768
rect 18748 17756 18754 17808
rect 27430 17756 27436 17808
rect 27488 17756 27494 17808
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 12032 17700 12265 17728
rect 12032 17688 12038 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 12345 17731 12403 17737
rect 12345 17697 12357 17731
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 16393 17731 16451 17737
rect 16393 17697 16405 17731
rect 16439 17728 16451 17731
rect 17310 17728 17316 17740
rect 16439 17700 17316 17728
rect 16439 17697 16451 17700
rect 16393 17691 16451 17697
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 10980 17592 11008 17620
rect 10704 17564 11008 17592
rect 11057 17595 11115 17601
rect 10505 17555 10563 17561
rect 10796 17536 10824 17564
rect 11057 17561 11069 17595
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 11425 17595 11483 17601
rect 11425 17561 11437 17595
rect 11471 17592 11483 17595
rect 12066 17592 12072 17604
rect 11471 17564 12072 17592
rect 11471 17561 11483 17564
rect 11425 17555 11483 17561
rect 8444 17496 8524 17524
rect 8444 17484 8450 17496
rect 9122 17484 9128 17536
rect 9180 17484 9186 17536
rect 10778 17484 10784 17536
rect 10836 17484 10842 17536
rect 10965 17527 11023 17533
rect 10965 17493 10977 17527
rect 11011 17524 11023 17527
rect 11072 17524 11100 17555
rect 12066 17552 12072 17564
rect 12124 17552 12130 17604
rect 12250 17552 12256 17604
rect 12308 17592 12314 17604
rect 12360 17592 12388 17691
rect 17310 17688 17316 17700
rect 17368 17688 17374 17740
rect 19245 17731 19303 17737
rect 19245 17697 19257 17731
rect 19291 17728 19303 17731
rect 19426 17728 19432 17740
rect 19291 17700 19432 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 19426 17688 19432 17700
rect 19484 17728 19490 17740
rect 20254 17728 20260 17740
rect 19484 17700 20260 17728
rect 19484 17688 19490 17700
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 21269 17731 21327 17737
rect 21269 17697 21281 17731
rect 21315 17728 21327 17731
rect 22094 17728 22100 17740
rect 21315 17700 22100 17728
rect 21315 17697 21327 17700
rect 21269 17691 21327 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 25225 17731 25283 17737
rect 25225 17697 25237 17731
rect 25271 17728 25283 17731
rect 27614 17728 27620 17740
rect 25271 17700 27620 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 16669 17663 16727 17669
rect 16669 17629 16681 17663
rect 16715 17660 16727 17663
rect 18414 17660 18420 17672
rect 16715 17632 18420 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 18414 17620 18420 17632
rect 18472 17620 18478 17672
rect 21634 17620 21640 17672
rect 21692 17660 21698 17672
rect 21818 17660 21824 17672
rect 21692 17632 21824 17660
rect 21692 17620 21698 17632
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 21913 17663 21971 17669
rect 21913 17629 21925 17663
rect 21959 17629 21971 17663
rect 21913 17623 21971 17629
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24670 17660 24676 17672
rect 24627 17632 24676 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 12802 17592 12808 17604
rect 12308 17564 12808 17592
rect 12308 17552 12314 17564
rect 12802 17552 12808 17564
rect 12860 17552 12866 17604
rect 15841 17595 15899 17601
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 16393 17595 16451 17601
rect 16393 17592 16405 17595
rect 15887 17564 16405 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 16393 17561 16405 17564
rect 16439 17561 16451 17595
rect 16393 17555 16451 17561
rect 19978 17552 19984 17604
rect 20036 17552 20042 17604
rect 20993 17595 21051 17601
rect 20993 17561 21005 17595
rect 21039 17561 21051 17595
rect 20993 17555 21051 17561
rect 11011 17496 11100 17524
rect 11011 17493 11023 17496
rect 10965 17487 11023 17493
rect 11698 17484 11704 17536
rect 11756 17524 11762 17536
rect 12161 17527 12219 17533
rect 12161 17524 12173 17527
rect 11756 17496 12173 17524
rect 11756 17484 11762 17496
rect 12161 17493 12173 17496
rect 12207 17493 12219 17527
rect 12161 17487 12219 17493
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 15102 17524 15108 17536
rect 12400 17496 15108 17524
rect 12400 17484 12406 17496
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 15344 17496 15485 17524
rect 15344 17484 15350 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 19702 17484 19708 17536
rect 19760 17524 19766 17536
rect 21008 17524 21036 17555
rect 19760 17496 21036 17524
rect 19760 17484 19766 17496
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 21929 17524 21957 17623
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 28905 17663 28963 17669
rect 28905 17660 28917 17663
rect 27580 17632 28917 17660
rect 27580 17620 27586 17632
rect 28905 17629 28917 17632
rect 28951 17629 28963 17663
rect 28905 17623 28963 17629
rect 25498 17552 25504 17604
rect 25556 17552 25562 17604
rect 26234 17552 26240 17604
rect 26292 17552 26298 17604
rect 26786 17552 26792 17604
rect 26844 17592 26850 17604
rect 27065 17595 27123 17601
rect 27065 17592 27077 17595
rect 26844 17564 27077 17592
rect 26844 17552 26850 17564
rect 27065 17561 27077 17564
rect 27111 17561 27123 17595
rect 27065 17555 27123 17561
rect 22094 17524 22100 17536
rect 21324 17496 22100 17524
rect 21324 17484 21330 17496
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 26326 17484 26332 17536
rect 26384 17524 26390 17536
rect 26973 17527 27031 17533
rect 26973 17524 26985 17527
rect 26384 17496 26985 17524
rect 26384 17484 26390 17496
rect 26973 17493 26985 17496
rect 27019 17524 27031 17527
rect 27154 17524 27160 17536
rect 27019 17496 27160 17524
rect 27019 17493 27031 17496
rect 26973 17487 27031 17493
rect 27154 17484 27160 17496
rect 27212 17484 27218 17536
rect 27525 17527 27583 17533
rect 27525 17493 27537 17527
rect 27571 17524 27583 17527
rect 27706 17524 27712 17536
rect 27571 17496 27712 17524
rect 27571 17493 27583 17496
rect 27525 17487 27583 17493
rect 27706 17484 27712 17496
rect 27764 17484 27770 17536
rect 1104 17434 29716 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 29716 17434
rect 1104 17360 29716 17382
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 3421 17323 3479 17329
rect 3421 17320 3433 17323
rect 3384 17292 3433 17320
rect 3384 17280 3390 17292
rect 3421 17289 3433 17292
rect 3467 17289 3479 17323
rect 3976 17323 4034 17329
rect 3976 17320 3988 17323
rect 3421 17283 3479 17289
rect 3896 17292 3988 17320
rect 842 17212 848 17264
rect 900 17252 906 17264
rect 1489 17255 1547 17261
rect 1489 17252 1501 17255
rect 900 17224 1501 17252
rect 900 17212 906 17224
rect 1489 17221 1501 17224
rect 1535 17221 1547 17255
rect 3694 17252 3700 17264
rect 1489 17215 1547 17221
rect 3436 17224 3700 17252
rect 3436 17193 3464 17224
rect 3694 17212 3700 17224
rect 3752 17252 3758 17264
rect 3896 17252 3924 17292
rect 3976 17289 3988 17292
rect 4022 17289 4034 17323
rect 3976 17283 4034 17289
rect 4249 17323 4307 17329
rect 4249 17289 4261 17323
rect 4295 17320 4307 17323
rect 4522 17320 4528 17332
rect 4295 17292 4528 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 5718 17320 5724 17332
rect 4632 17292 5724 17320
rect 4632 17252 4660 17292
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 6914 17280 6920 17332
rect 6972 17280 6978 17332
rect 7098 17280 7104 17332
rect 7156 17280 7162 17332
rect 7558 17320 7564 17332
rect 7392 17292 7564 17320
rect 7392 17252 7420 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 10226 17320 10232 17332
rect 7708 17292 10232 17320
rect 7708 17280 7714 17292
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 10410 17280 10416 17332
rect 10468 17320 10474 17332
rect 10962 17320 10968 17332
rect 10468 17292 10968 17320
rect 10468 17280 10474 17292
rect 10962 17280 10968 17292
rect 11020 17280 11026 17332
rect 18601 17323 18659 17329
rect 18601 17289 18613 17323
rect 18647 17320 18659 17323
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 18647 17292 19349 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 19702 17280 19708 17332
rect 19760 17280 19766 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 20073 17323 20131 17329
rect 20073 17320 20085 17323
rect 20036 17292 20085 17320
rect 20036 17280 20042 17292
rect 20073 17289 20085 17292
rect 20119 17289 20131 17323
rect 20073 17283 20131 17289
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 21416 17292 21496 17320
rect 21416 17280 21422 17292
rect 3752 17224 3924 17252
rect 4448 17224 4660 17252
rect 4724 17224 7420 17252
rect 7469 17255 7527 17261
rect 3752 17212 3758 17224
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17153 3663 17187
rect 3605 17147 3663 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 3620 17116 3648 17147
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 3881 17187 3939 17193
rect 3881 17153 3893 17187
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 4338 17184 4344 17196
rect 4295 17156 4344 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 3896 17116 3924 17147
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 4448 17193 4476 17224
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 4617 17190 4675 17193
rect 4724 17190 4752 17224
rect 7469 17221 7481 17255
rect 7515 17252 7527 17255
rect 10321 17255 10379 17261
rect 7515 17224 8800 17252
rect 7515 17221 7527 17224
rect 7469 17215 7527 17221
rect 4617 17187 4752 17190
rect 4617 17153 4629 17187
rect 4663 17162 4752 17187
rect 4663 17153 4675 17162
rect 4617 17147 4675 17153
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 8294 17184 8300 17196
rect 7607 17156 8300 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 4706 17116 4712 17128
rect 1719 17088 2774 17116
rect 3620 17088 4712 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2746 16980 2774 17088
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7650 17076 7656 17128
rect 7708 17076 7714 17128
rect 8386 17076 8392 17128
rect 8444 17076 8450 17128
rect 8772 17125 8800 17224
rect 10321 17221 10333 17255
rect 10367 17252 10379 17255
rect 11241 17255 11299 17261
rect 11241 17252 11253 17255
rect 10367 17224 11253 17252
rect 10367 17221 10379 17224
rect 10321 17215 10379 17221
rect 11241 17221 11253 17224
rect 11287 17221 11299 17255
rect 11241 17215 11299 17221
rect 12360 17224 13308 17252
rect 9125 17187 9183 17193
rect 9125 17153 9137 17187
rect 9171 17184 9183 17187
rect 9674 17184 9680 17196
rect 9171 17156 9680 17184
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17085 8815 17119
rect 8757 17079 8815 17085
rect 4111 17051 4169 17057
rect 4111 17017 4123 17051
rect 4157 17048 4169 17051
rect 4433 17051 4491 17057
rect 4433 17048 4445 17051
rect 4157 17020 4445 17048
rect 4157 17017 4169 17020
rect 4111 17011 4169 17017
rect 4433 17017 4445 17020
rect 4479 17017 4491 17051
rect 4433 17011 4491 17017
rect 4614 17008 4620 17060
rect 4672 17048 4678 17060
rect 7834 17048 7840 17060
rect 4672 17020 7840 17048
rect 4672 17008 4678 17020
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 8665 17051 8723 17057
rect 8665 17017 8677 17051
rect 8711 17048 8723 17051
rect 9140 17048 9168 17147
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10594 17193 10600 17196
rect 10551 17187 10600 17193
rect 10551 17153 10563 17187
rect 10597 17153 10600 17187
rect 10551 17147 10600 17153
rect 10594 17144 10600 17147
rect 10652 17144 10658 17196
rect 10686 17144 10692 17196
rect 10744 17144 10750 17196
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17116 9275 17119
rect 10045 17119 10103 17125
rect 10045 17116 10057 17119
rect 9263 17088 10057 17116
rect 9263 17085 9275 17088
rect 9217 17079 9275 17085
rect 10045 17085 10057 17088
rect 10091 17085 10103 17119
rect 10244 17116 10272 17144
rect 10796 17116 10824 17147
rect 10962 17144 10968 17196
rect 11020 17144 11026 17196
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 12360 17193 12388 17224
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 11388 17156 12357 17184
rect 11388 17144 11394 17156
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 12345 17147 12403 17153
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 10244 17088 10824 17116
rect 10873 17119 10931 17125
rect 10045 17079 10103 17085
rect 10873 17085 10885 17119
rect 10919 17116 10931 17119
rect 12544 17116 12572 17147
rect 12802 17144 12808 17196
rect 12860 17144 12866 17196
rect 13280 17193 13308 17224
rect 16224 17224 18368 17252
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17184 13323 17187
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13311 17156 13461 17184
rect 13311 17153 13323 17156
rect 13265 17147 13323 17153
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 13096 17116 13124 17147
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 16224 17193 16252 17224
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13780 17156 14105 17184
rect 13780 17144 13786 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 10919 17088 13124 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 13998 17076 14004 17128
rect 14056 17076 14062 17128
rect 14274 17076 14280 17128
rect 14332 17116 14338 17128
rect 15010 17116 15016 17128
rect 14332 17088 15016 17116
rect 14332 17076 14338 17088
rect 15010 17076 15016 17088
rect 15068 17116 15074 17128
rect 16224 17116 16252 17147
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 18340 17184 18368 17224
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 19242 17252 19248 17264
rect 18472 17224 19248 17252
rect 18472 17212 18478 17224
rect 19242 17212 19248 17224
rect 19300 17252 19306 17264
rect 21468 17261 21496 17292
rect 21542 17280 21548 17332
rect 21600 17320 21606 17332
rect 21600 17292 21864 17320
rect 21600 17280 21606 17292
rect 20533 17255 20591 17261
rect 20533 17252 20545 17255
rect 19300 17224 20545 17252
rect 19300 17212 19306 17224
rect 20533 17221 20545 17224
rect 20579 17221 20591 17255
rect 20533 17215 20591 17221
rect 21453 17255 21511 17261
rect 21453 17221 21465 17255
rect 21499 17252 21511 17255
rect 21726 17252 21732 17264
rect 21499 17224 21732 17252
rect 21499 17221 21511 17224
rect 21453 17215 21511 17221
rect 21726 17212 21732 17224
rect 21784 17212 21790 17264
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 18340 17156 19993 17184
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17184 20683 17187
rect 21358 17184 21364 17196
rect 20671 17156 21364 17184
rect 20671 17153 20683 17156
rect 20625 17147 20683 17153
rect 21358 17144 21364 17156
rect 21416 17144 21422 17196
rect 21634 17144 21640 17196
rect 21692 17144 21698 17196
rect 21836 17193 21864 17292
rect 22094 17280 22100 17332
rect 22152 17280 22158 17332
rect 26513 17323 26571 17329
rect 26513 17289 26525 17323
rect 26559 17320 26571 17323
rect 27062 17320 27068 17332
rect 26559 17292 27068 17320
rect 26559 17289 26571 17292
rect 26513 17283 26571 17289
rect 27062 17280 27068 17292
rect 27120 17320 27126 17332
rect 29181 17323 29239 17329
rect 29181 17320 29193 17323
rect 27120 17292 29193 17320
rect 27120 17280 27126 17292
rect 29181 17289 29193 17292
rect 29227 17289 29239 17323
rect 29181 17283 29239 17289
rect 22112 17252 22140 17280
rect 26421 17255 26479 17261
rect 26421 17252 26433 17255
rect 22112 17224 22329 17252
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 15068 17088 16252 17116
rect 15068 17076 15074 17088
rect 18138 17076 18144 17128
rect 18196 17076 18202 17128
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 19245 17119 19303 17125
rect 19245 17085 19257 17119
rect 19291 17116 19303 17119
rect 19426 17116 19432 17128
rect 19291 17088 19432 17116
rect 19291 17085 19303 17088
rect 19245 17079 19303 17085
rect 8711 17020 9168 17048
rect 8711 17017 8723 17020
rect 8665 17011 8723 17017
rect 12894 17008 12900 17060
rect 12952 17048 12958 17060
rect 13173 17051 13231 17057
rect 13173 17048 13185 17051
rect 12952 17020 13185 17048
rect 12952 17008 12958 17020
rect 13173 17017 13185 17020
rect 13219 17017 13231 17051
rect 19168 17048 19196 17079
rect 19426 17076 19432 17088
rect 19484 17076 19490 17128
rect 21836 17116 21864 17147
rect 21910 17144 21916 17196
rect 21968 17184 21974 17196
rect 21968 17156 22013 17184
rect 21968 17144 21974 17156
rect 22094 17144 22100 17196
rect 22152 17144 22158 17196
rect 22301 17193 22329 17224
rect 25608 17224 26433 17252
rect 25608 17196 25636 17224
rect 26421 17221 26433 17224
rect 26467 17221 26479 17255
rect 26421 17215 26479 17221
rect 26786 17212 26792 17264
rect 26844 17212 26850 17264
rect 27614 17252 27620 17264
rect 27448 17224 27620 17252
rect 22189 17187 22247 17193
rect 22189 17153 22201 17187
rect 22235 17153 22247 17187
rect 22189 17147 22247 17153
rect 22286 17187 22344 17193
rect 22286 17153 22298 17187
rect 22332 17153 22344 17187
rect 22286 17147 22344 17153
rect 19812 17088 21864 17116
rect 19812 17060 19840 17088
rect 19794 17048 19800 17060
rect 19168 17020 19800 17048
rect 13173 17011 13231 17017
rect 19794 17008 19800 17020
rect 19852 17008 19858 17060
rect 12342 16980 12348 16992
rect 2746 16952 12348 16980
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 12989 16983 13047 16989
rect 12989 16980 13001 16983
rect 12768 16952 13001 16980
rect 12768 16940 12774 16952
rect 12989 16949 13001 16952
rect 13035 16949 13047 16983
rect 12989 16943 13047 16949
rect 16301 16983 16359 16989
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 16574 16980 16580 16992
rect 16347 16952 16580 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21634 16980 21640 16992
rect 21315 16952 21640 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21634 16940 21640 16952
rect 21692 16980 21698 16992
rect 22204 16980 22232 17147
rect 25590 17144 25596 17196
rect 25648 17144 25654 17196
rect 25777 17187 25835 17193
rect 25777 17153 25789 17187
rect 25823 17153 25835 17187
rect 25777 17147 25835 17153
rect 26237 17187 26295 17193
rect 26237 17153 26249 17187
rect 26283 17184 26295 17187
rect 26326 17184 26332 17196
rect 26283 17156 26332 17184
rect 26283 17153 26295 17156
rect 26237 17147 26295 17153
rect 25792 17116 25820 17147
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 27448 17193 27476 17224
rect 27614 17212 27620 17224
rect 27672 17212 27678 17264
rect 27706 17212 27712 17264
rect 27764 17212 27770 17264
rect 28718 17212 28724 17264
rect 28776 17212 28782 17264
rect 26605 17187 26663 17193
rect 26605 17153 26617 17187
rect 26651 17153 26663 17187
rect 26605 17147 26663 17153
rect 27433 17187 27491 17193
rect 27433 17153 27445 17187
rect 27479 17153 27491 17187
rect 27433 17147 27491 17153
rect 26050 17116 26056 17128
rect 25792 17088 26056 17116
rect 26050 17076 26056 17088
rect 26108 17116 26114 17128
rect 26620 17116 26648 17147
rect 26108 17088 26648 17116
rect 26108 17076 26114 17088
rect 21692 16952 22232 16980
rect 21692 16940 21698 16952
rect 22370 16940 22376 16992
rect 22428 16980 22434 16992
rect 22465 16983 22523 16989
rect 22465 16980 22477 16983
rect 22428 16952 22477 16980
rect 22428 16940 22434 16952
rect 22465 16949 22477 16952
rect 22511 16949 22523 16983
rect 22465 16943 22523 16949
rect 25406 16940 25412 16992
rect 25464 16940 25470 16992
rect 1104 16890 29716 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 29716 16890
rect 1104 16816 29716 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 17954 16776 17960 16788
rect 1627 16748 17960 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18138 16736 18144 16788
rect 18196 16736 18202 16788
rect 20898 16736 20904 16788
rect 20956 16736 20962 16788
rect 21177 16779 21235 16785
rect 21177 16745 21189 16779
rect 21223 16776 21235 16779
rect 21266 16776 21272 16788
rect 21223 16748 21272 16776
rect 21223 16745 21235 16748
rect 21177 16739 21235 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 21453 16779 21511 16785
rect 21453 16745 21465 16779
rect 21499 16745 21511 16779
rect 25590 16776 25596 16788
rect 21453 16739 21511 16745
rect 25056 16748 25596 16776
rect 5718 16668 5724 16720
rect 5776 16708 5782 16720
rect 8386 16708 8392 16720
rect 5776 16680 8392 16708
rect 5776 16668 5782 16680
rect 2866 16600 2872 16652
rect 2924 16640 2930 16652
rect 6822 16640 6828 16652
rect 2924 16612 6828 16640
rect 2924 16600 2930 16612
rect 842 16532 848 16584
rect 900 16572 906 16584
rect 6564 16581 6592 16612
rect 6822 16600 6828 16612
rect 6880 16600 6886 16652
rect 7576 16649 7604 16680
rect 8386 16668 8392 16680
rect 8444 16668 8450 16720
rect 14642 16708 14648 16720
rect 10428 16680 14648 16708
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8846 16640 8852 16652
rect 7883 16612 8852 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 10318 16640 10324 16652
rect 10244 16612 10324 16640
rect 1489 16575 1547 16581
rect 1489 16572 1501 16575
rect 900 16544 1501 16572
rect 900 16532 906 16544
rect 1489 16541 1501 16544
rect 1535 16541 1547 16575
rect 1489 16535 1547 16541
rect 6549 16575 6607 16581
rect 6549 16541 6561 16575
rect 6595 16541 6607 16575
rect 6549 16535 6607 16541
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 7340 16544 7481 16572
rect 7340 16532 7346 16544
rect 7469 16541 7481 16544
rect 7515 16572 7527 16575
rect 8202 16572 8208 16584
rect 7515 16544 8208 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 8202 16532 8208 16544
rect 8260 16572 8266 16584
rect 9858 16572 9864 16584
rect 8260 16544 9864 16572
rect 8260 16532 8266 16544
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 10244 16581 10272 16612
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10428 16581 10456 16680
rect 14642 16668 14648 16680
rect 14700 16668 14706 16720
rect 17402 16668 17408 16720
rect 17460 16708 17466 16720
rect 18046 16708 18052 16720
rect 17460 16680 18052 16708
rect 17460 16668 17466 16680
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 21468 16708 21496 16739
rect 21192 16680 21496 16708
rect 22833 16711 22891 16717
rect 21192 16652 21220 16680
rect 22833 16677 22845 16711
rect 22879 16708 22891 16711
rect 24486 16708 24492 16720
rect 22879 16680 24492 16708
rect 22879 16677 22891 16680
rect 22833 16671 22891 16677
rect 24486 16668 24492 16680
rect 24544 16668 24550 16720
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 15197 16643 15255 16649
rect 15197 16640 15209 16643
rect 13504 16612 15209 16640
rect 13504 16600 13510 16612
rect 15197 16609 15209 16612
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 16666 16600 16672 16652
rect 16724 16640 16730 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16724 16612 17233 16640
rect 16724 16600 16730 16612
rect 17221 16609 17233 16612
rect 17267 16640 17279 16643
rect 17267 16612 18460 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10413 16575 10471 16581
rect 10413 16541 10425 16575
rect 10459 16541 10471 16575
rect 10413 16535 10471 16541
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16541 10655 16575
rect 10597 16535 10655 16541
rect 10751 16575 10809 16581
rect 10751 16541 10763 16575
rect 10797 16572 10809 16575
rect 10962 16572 10968 16584
rect 10797 16544 10968 16572
rect 10797 16541 10809 16544
rect 10751 16535 10809 16541
rect 1578 16464 1584 16516
rect 1636 16504 1642 16516
rect 7006 16504 7012 16516
rect 1636 16476 7012 16504
rect 1636 16464 1642 16476
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 10612 16504 10640 16535
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 12710 16532 12716 16584
rect 12768 16532 12774 16584
rect 12894 16532 12900 16584
rect 12952 16532 12958 16584
rect 13078 16532 13084 16584
rect 13136 16532 13142 16584
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 16574 16532 16580 16584
rect 16632 16532 16638 16584
rect 17402 16532 17408 16584
rect 17460 16532 17466 16584
rect 17595 16581 17623 16612
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 17675 16575 17733 16581
rect 17675 16541 17687 16575
rect 17721 16541 17733 16575
rect 17675 16535 17733 16541
rect 17773 16575 17831 16581
rect 17773 16541 17785 16575
rect 17819 16572 17831 16575
rect 17862 16572 17868 16584
rect 17819 16544 17868 16572
rect 17819 16541 17831 16544
rect 17773 16535 17831 16541
rect 10336 16476 10640 16504
rect 12989 16507 13047 16513
rect 6638 16396 6644 16448
rect 6696 16396 6702 16448
rect 10042 16396 10048 16448
rect 10100 16436 10106 16448
rect 10336 16445 10364 16476
rect 12989 16473 13001 16507
rect 13035 16504 13047 16507
rect 13722 16504 13728 16516
rect 13035 16476 13728 16504
rect 13035 16473 13047 16476
rect 12989 16467 13047 16473
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 15470 16464 15476 16516
rect 15528 16464 15534 16516
rect 17696 16504 17724 16535
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 17954 16532 17960 16584
rect 18012 16532 18018 16584
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18432 16581 18460 16612
rect 20254 16600 20260 16652
rect 20312 16640 20318 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20312 16612 20821 16640
rect 20312 16600 20318 16612
rect 20809 16609 20821 16612
rect 20855 16609 20867 16643
rect 20809 16603 20867 16609
rect 21174 16600 21180 16652
rect 21232 16600 21238 16652
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 21545 16643 21603 16649
rect 21545 16640 21557 16643
rect 21416 16612 21557 16640
rect 21416 16600 21422 16612
rect 21545 16609 21557 16612
rect 21591 16640 21603 16643
rect 21591 16612 22094 16640
rect 21591 16609 21603 16612
rect 21545 16603 21603 16609
rect 18233 16575 18291 16581
rect 18233 16572 18245 16575
rect 18104 16544 18245 16572
rect 18104 16532 18110 16544
rect 18233 16541 18245 16544
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 19702 16572 19708 16584
rect 18463 16544 19708 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 21634 16532 21640 16584
rect 21692 16532 21698 16584
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 17696 16476 17816 16504
rect 17788 16448 17816 16476
rect 20346 16464 20352 16516
rect 20404 16504 20410 16516
rect 20717 16507 20775 16513
rect 20717 16504 20729 16507
rect 20404 16476 20729 16504
rect 20404 16464 20410 16476
rect 20717 16473 20729 16476
rect 20763 16473 20775 16507
rect 20717 16467 20775 16473
rect 21542 16464 21548 16516
rect 21600 16504 21606 16516
rect 21744 16504 21772 16535
rect 21818 16532 21824 16584
rect 21876 16572 21882 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21876 16544 21925 16572
rect 21876 16532 21882 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 22066 16572 22094 16612
rect 22370 16600 22376 16652
rect 22428 16600 22434 16652
rect 22462 16572 22468 16584
rect 22066 16544 22468 16572
rect 21913 16535 21971 16541
rect 22462 16532 22468 16544
rect 22520 16532 22526 16584
rect 24213 16575 24271 16581
rect 24213 16541 24225 16575
rect 24259 16572 24271 16575
rect 24670 16572 24676 16584
rect 24259 16544 24676 16572
rect 24259 16541 24271 16544
rect 24213 16535 24271 16541
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 25056 16581 25084 16748
rect 25590 16736 25596 16748
rect 25648 16776 25654 16788
rect 26881 16779 26939 16785
rect 26881 16776 26893 16779
rect 25648 16748 26893 16776
rect 25648 16736 25654 16748
rect 26881 16745 26893 16748
rect 26927 16745 26939 16779
rect 26881 16739 26939 16745
rect 26896 16708 26924 16739
rect 27430 16736 27436 16788
rect 27488 16776 27494 16788
rect 27525 16779 27583 16785
rect 27525 16776 27537 16779
rect 27488 16748 27537 16776
rect 27488 16736 27494 16748
rect 27525 16745 27537 16748
rect 27571 16745 27583 16779
rect 27525 16739 27583 16745
rect 28629 16779 28687 16785
rect 28629 16745 28641 16779
rect 28675 16776 28687 16779
rect 28718 16776 28724 16788
rect 28675 16748 28724 16776
rect 28675 16745 28687 16748
rect 28629 16739 28687 16745
rect 28718 16736 28724 16748
rect 28776 16736 28782 16788
rect 26896 16680 27292 16708
rect 25130 16600 25136 16652
rect 25188 16600 25194 16652
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 26108 16612 27016 16640
rect 26108 16600 26114 16612
rect 24857 16575 24915 16581
rect 24857 16541 24869 16575
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 25041 16575 25099 16581
rect 25041 16541 25053 16575
rect 25087 16541 25099 16575
rect 26988 16572 27016 16612
rect 27062 16600 27068 16652
rect 27120 16600 27126 16652
rect 27154 16600 27160 16652
rect 27212 16600 27218 16652
rect 27264 16649 27292 16680
rect 29086 16668 29092 16720
rect 29144 16668 29150 16720
rect 27249 16643 27307 16649
rect 27249 16609 27261 16643
rect 27295 16609 27307 16643
rect 27249 16603 27307 16609
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16609 27399 16643
rect 27341 16603 27399 16609
rect 27356 16572 27384 16603
rect 27430 16600 27436 16652
rect 27488 16640 27494 16652
rect 27488 16612 29040 16640
rect 27488 16600 27494 16612
rect 26988 16544 27384 16572
rect 25041 16535 25099 16541
rect 21600 16476 21772 16504
rect 24872 16504 24900 16535
rect 28166 16532 28172 16584
rect 28224 16572 28230 16584
rect 28736 16581 28764 16612
rect 29012 16581 29040 16612
rect 28261 16575 28319 16581
rect 28261 16572 28273 16575
rect 28224 16544 28273 16572
rect 28224 16532 28230 16544
rect 28261 16541 28273 16544
rect 28307 16541 28319 16575
rect 28261 16535 28319 16541
rect 28721 16575 28779 16581
rect 28721 16541 28733 16575
rect 28767 16541 28779 16575
rect 28721 16535 28779 16541
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 29270 16532 29276 16584
rect 29328 16532 29334 16584
rect 25409 16507 25467 16513
rect 24872 16476 25176 16504
rect 21600 16464 21606 16476
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 10100 16408 10333 16436
rect 10100 16396 10106 16408
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 10321 16399 10379 16405
rect 10962 16396 10968 16448
rect 11020 16396 11026 16448
rect 13265 16439 13323 16445
rect 13265 16405 13277 16439
rect 13311 16436 13323 16439
rect 13538 16436 13544 16448
rect 13311 16408 13544 16436
rect 13311 16405 13323 16408
rect 13265 16399 13323 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14332 16408 14381 16436
rect 14332 16396 14338 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14369 16399 14427 16405
rect 17494 16396 17500 16448
rect 17552 16396 17558 16448
rect 17770 16396 17776 16448
rect 17828 16396 17834 16448
rect 17862 16396 17868 16448
rect 17920 16436 17926 16448
rect 18325 16439 18383 16445
rect 18325 16436 18337 16439
rect 17920 16408 18337 16436
rect 17920 16396 17926 16408
rect 18325 16405 18337 16408
rect 18371 16405 18383 16439
rect 18325 16399 18383 16405
rect 21266 16396 21272 16448
rect 21324 16396 21330 16448
rect 21913 16439 21971 16445
rect 21913 16405 21925 16439
rect 21959 16436 21971 16439
rect 22094 16436 22100 16448
rect 21959 16408 22100 16436
rect 21959 16405 21971 16408
rect 21913 16399 21971 16405
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 24121 16439 24179 16445
rect 24121 16436 24133 16439
rect 24084 16408 24133 16436
rect 24084 16396 24090 16408
rect 24121 16405 24133 16408
rect 24167 16405 24179 16439
rect 24121 16399 24179 16405
rect 25038 16396 25044 16448
rect 25096 16396 25102 16448
rect 25148 16436 25176 16476
rect 25409 16473 25421 16507
rect 25455 16504 25467 16507
rect 25498 16504 25504 16516
rect 25455 16476 25504 16504
rect 25455 16473 25467 16476
rect 25409 16467 25467 16473
rect 25498 16464 25504 16476
rect 25556 16464 25562 16516
rect 26418 16464 26424 16516
rect 26476 16464 26482 16516
rect 26050 16436 26056 16448
rect 25148 16408 26056 16436
rect 26050 16396 26056 16408
rect 26108 16396 26114 16448
rect 28442 16396 28448 16448
rect 28500 16396 28506 16448
rect 28902 16396 28908 16448
rect 28960 16396 28966 16448
rect 1104 16346 29716 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 29716 16346
rect 1104 16272 29716 16294
rect 5994 16232 6000 16244
rect 1688 16204 6000 16232
rect 1688 16105 1716 16204
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6564 16204 9076 16232
rect 2590 16124 2596 16176
rect 2648 16124 2654 16176
rect 3697 16167 3755 16173
rect 3697 16133 3709 16167
rect 3743 16164 3755 16167
rect 3786 16164 3792 16176
rect 3743 16136 3792 16164
rect 3743 16133 3755 16136
rect 3697 16127 3755 16133
rect 3786 16124 3792 16136
rect 3844 16164 3850 16176
rect 4157 16167 4215 16173
rect 3844 16136 4108 16164
rect 3844 16124 3850 16136
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 3326 16056 3332 16108
rect 3384 16096 3390 16108
rect 3878 16096 3884 16108
rect 3384 16068 3884 16096
rect 3384 16056 3390 16068
rect 3878 16056 3884 16068
rect 3936 16096 3942 16108
rect 4080 16105 4108 16136
rect 4157 16133 4169 16167
rect 4203 16164 4215 16167
rect 4706 16164 4712 16176
rect 4203 16136 4712 16164
rect 4203 16133 4215 16136
rect 4157 16127 4215 16133
rect 4706 16124 4712 16136
rect 4764 16164 4770 16176
rect 5442 16164 5448 16176
rect 4764 16136 5448 16164
rect 4764 16124 4770 16136
rect 5442 16124 5448 16136
rect 5500 16124 5506 16176
rect 5537 16167 5595 16173
rect 5537 16133 5549 16167
rect 5583 16164 5595 16167
rect 6564 16164 6592 16204
rect 9048 16176 9076 16204
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9217 16235 9275 16241
rect 9217 16232 9229 16235
rect 9180 16204 9229 16232
rect 9180 16192 9186 16204
rect 9217 16201 9229 16204
rect 9263 16201 9275 16235
rect 9217 16195 9275 16201
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10505 16235 10563 16241
rect 10505 16232 10517 16235
rect 10376 16204 10517 16232
rect 10376 16192 10382 16204
rect 10505 16201 10517 16204
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11698 16232 11704 16244
rect 11379 16204 11704 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 12124 16204 12173 16232
rect 12124 16192 12130 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 13780 16204 14872 16232
rect 13780 16192 13786 16204
rect 5583 16136 6592 16164
rect 5583 16133 5595 16136
rect 5537 16127 5595 16133
rect 6638 16124 6644 16176
rect 6696 16164 6702 16176
rect 6696 16136 7130 16164
rect 6696 16124 6702 16136
rect 8202 16124 8208 16176
rect 8260 16164 8266 16176
rect 8389 16167 8447 16173
rect 8389 16164 8401 16167
rect 8260 16136 8401 16164
rect 8260 16124 8266 16136
rect 8389 16133 8401 16136
rect 8435 16133 8447 16167
rect 8389 16127 8447 16133
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 9088 16136 11744 16164
rect 9088 16124 9094 16136
rect 3973 16099 4031 16105
rect 3973 16096 3985 16099
rect 3936 16068 3985 16096
rect 3936 16056 3942 16068
rect 3973 16065 3985 16068
rect 4019 16065 4031 16099
rect 3973 16059 4031 16065
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 4111 16094 4200 16096
rect 4246 16094 4252 16108
rect 4111 16068 4252 16094
rect 4111 16065 4123 16068
rect 4172 16066 4252 16068
rect 4065 16059 4123 16065
rect 4246 16056 4252 16066
rect 4304 16056 4310 16108
rect 4341 16099 4399 16105
rect 4341 16065 4353 16099
rect 4387 16065 4399 16099
rect 4341 16059 4399 16065
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 1995 16000 3280 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 3252 15960 3280 16000
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 4356 16028 4384 16059
rect 4614 16056 4620 16108
rect 4672 16056 4678 16108
rect 4801 16099 4859 16105
rect 4801 16065 4813 16099
rect 4847 16096 4859 16099
rect 4847 16068 5120 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 3660 16000 4384 16028
rect 3660 15988 3666 16000
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 3252 15932 3801 15960
rect 3789 15929 3801 15932
rect 3835 15929 3847 15963
rect 3789 15923 3847 15929
rect 3970 15920 3976 15972
rect 4028 15960 4034 15972
rect 5092 15960 5120 16068
rect 5166 16056 5172 16108
rect 5224 16056 5230 16108
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5276 16028 5304 16059
rect 5350 16056 5356 16108
rect 5408 16056 5414 16108
rect 5994 16056 6000 16108
rect 6052 16096 6058 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6052 16068 6377 16096
rect 6052 16056 6058 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 8846 16056 8852 16108
rect 8904 16096 8910 16108
rect 9140 16105 9168 16136
rect 9125 16099 9183 16105
rect 8904 16068 9076 16096
rect 8904 16056 8910 16068
rect 5626 16028 5632 16040
rect 5276 16000 5632 16028
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 6638 15988 6644 16040
rect 6696 15988 6702 16040
rect 8938 15988 8944 16040
rect 8996 15988 9002 16040
rect 9048 16028 9076 16068
rect 9125 16065 9137 16099
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 9674 16056 9680 16108
rect 9732 16056 9738 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 9048 16000 9597 16028
rect 9585 15997 9597 16000
rect 9631 16028 9643 16031
rect 9876 16028 9904 16059
rect 9631 16000 9904 16028
rect 9968 16028 9996 16059
rect 10042 16056 10048 16108
rect 10100 16056 10106 16108
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16065 10287 16099
rect 10229 16059 10287 16065
rect 10329 16099 10387 16105
rect 10329 16065 10341 16099
rect 10375 16096 10387 16099
rect 10778 16096 10784 16108
rect 10375 16068 10784 16096
rect 10375 16065 10387 16068
rect 10329 16059 10387 16065
rect 9968 16000 10088 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 10060 15972 10088 16000
rect 5718 15960 5724 15972
rect 4028 15932 5724 15960
rect 4028 15920 4034 15932
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 9401 15963 9459 15969
rect 9401 15929 9413 15963
rect 9447 15960 9459 15963
rect 10042 15960 10048 15972
rect 9447 15932 10048 15960
rect 9447 15929 9459 15932
rect 9401 15923 9459 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4614 15892 4620 15904
rect 4479 15864 4620 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 9766 15852 9772 15904
rect 9824 15852 9830 15904
rect 9858 15852 9864 15904
rect 9916 15892 9922 15904
rect 10244 15892 10272 16059
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 10428 15960 10456 16068
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10962 16056 10968 16108
rect 11020 16056 11026 16108
rect 11716 16105 11744 16136
rect 11790 16124 11796 16176
rect 11848 16164 11854 16176
rect 13446 16164 13452 16176
rect 11848 16136 13452 16164
rect 11848 16124 11854 16136
rect 13280 16105 13308 16136
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 13538 16124 13544 16176
rect 13596 16124 13602 16176
rect 14274 16124 14280 16176
rect 14332 16124 14338 16176
rect 14844 16164 14872 16204
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 15565 16235 15623 16241
rect 15565 16232 15577 16235
rect 15528 16204 15577 16232
rect 15528 16192 15534 16204
rect 15565 16201 15577 16204
rect 15611 16201 15623 16235
rect 15565 16195 15623 16201
rect 16025 16235 16083 16241
rect 16025 16201 16037 16235
rect 16071 16232 16083 16235
rect 16666 16232 16672 16244
rect 16071 16204 16672 16232
rect 16071 16201 16083 16204
rect 16025 16195 16083 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 19610 16232 19616 16244
rect 18748 16204 19616 16232
rect 18748 16192 18754 16204
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 20714 16232 20720 16244
rect 20211 16204 20720 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 20901 16235 20959 16241
rect 20901 16201 20913 16235
rect 20947 16232 20959 16235
rect 20947 16204 22094 16232
rect 20947 16201 20959 16204
rect 20901 16195 20959 16201
rect 15289 16167 15347 16173
rect 15289 16164 15301 16167
rect 14844 16136 15301 16164
rect 15289 16133 15301 16136
rect 15335 16133 15347 16167
rect 15289 16127 15347 16133
rect 17770 16124 17776 16176
rect 17828 16164 17834 16176
rect 17828 16136 20117 16164
rect 17828 16124 17834 16136
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 12164 16099 12222 16105
rect 12164 16065 12176 16099
rect 12210 16065 12222 16099
rect 12164 16059 12222 16065
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16065 13323 16099
rect 13265 16059 13323 16065
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 10873 16031 10931 16037
rect 10873 16028 10885 16031
rect 10560 16000 10885 16028
rect 10560 15988 10566 16000
rect 10873 15997 10885 16000
rect 10919 15997 10931 16031
rect 10873 15991 10931 15997
rect 12176 15960 12204 16059
rect 15930 16056 15936 16108
rect 15988 16056 15994 16108
rect 19153 16099 19211 16105
rect 19153 16065 19165 16099
rect 19199 16096 19211 16099
rect 19334 16096 19340 16108
rect 19199 16068 19340 16096
rect 19199 16065 19211 16068
rect 19153 16059 19211 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19702 16056 19708 16108
rect 19760 16056 19766 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19904 16068 19993 16096
rect 14274 15988 14280 16040
rect 14332 16028 14338 16040
rect 16114 16028 16120 16040
rect 14332 16000 16120 16028
rect 14332 15988 14338 16000
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17862 16028 17868 16040
rect 17644 16000 17868 16028
rect 17644 15988 17650 16000
rect 17862 15988 17868 16000
rect 17920 16028 17926 16040
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17920 16000 18061 16028
rect 17920 15988 17926 16000
rect 18049 15997 18061 16000
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 19061 16031 19119 16037
rect 19061 16028 19073 16031
rect 18196 16000 19073 16028
rect 18196 15988 18202 16000
rect 19061 15997 19073 16000
rect 19107 16028 19119 16031
rect 19242 16028 19248 16040
rect 19107 16000 19248 16028
rect 19107 15997 19119 16000
rect 19061 15991 19119 15997
rect 19242 15988 19248 16000
rect 19300 15988 19306 16040
rect 12894 15960 12900 15972
rect 10376 15932 12900 15960
rect 10376 15920 10382 15932
rect 12894 15920 12900 15932
rect 12952 15920 12958 15972
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 17681 15963 17739 15969
rect 17681 15960 17693 15963
rect 17552 15932 17693 15960
rect 17552 15920 17558 15932
rect 17681 15929 17693 15932
rect 17727 15960 17739 15963
rect 17954 15960 17960 15972
rect 17727 15932 17960 15960
rect 17727 15929 17739 15932
rect 17681 15923 17739 15929
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 18785 15963 18843 15969
rect 18785 15929 18797 15963
rect 18831 15960 18843 15963
rect 18874 15960 18880 15972
rect 18831 15932 18880 15960
rect 18831 15929 18843 15932
rect 18785 15923 18843 15929
rect 18874 15920 18880 15932
rect 18932 15920 18938 15972
rect 19352 15960 19380 16056
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19484 16000 19809 16028
rect 19484 15988 19490 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 19904 15960 19932 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 20089 16096 20117 16136
rect 20254 16105 20260 16108
rect 20245 16099 20260 16105
rect 20245 16096 20257 16099
rect 20089 16068 20257 16096
rect 19981 16059 20039 16065
rect 20245 16065 20257 16068
rect 20245 16059 20260 16065
rect 20254 16056 20260 16059
rect 20312 16056 20318 16108
rect 20346 16056 20352 16108
rect 20404 16056 20410 16108
rect 20776 16099 20834 16105
rect 20776 16065 20788 16099
rect 20822 16096 20834 16099
rect 20898 16096 20904 16108
rect 20822 16068 20904 16096
rect 20822 16065 20834 16068
rect 20776 16059 20834 16065
rect 20898 16056 20904 16068
rect 20956 16056 20962 16108
rect 22066 16096 22094 16204
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22520 16204 23029 16232
rect 22520 16192 22526 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 23017 16195 23075 16201
rect 24670 16192 24676 16244
rect 24728 16192 24734 16244
rect 25498 16192 25504 16244
rect 25556 16232 25562 16244
rect 25593 16235 25651 16241
rect 25593 16232 25605 16235
rect 25556 16204 25605 16232
rect 25556 16192 25562 16204
rect 25593 16201 25605 16204
rect 25639 16201 25651 16235
rect 25593 16195 25651 16201
rect 26237 16235 26295 16241
rect 26237 16201 26249 16235
rect 26283 16232 26295 16235
rect 26418 16232 26424 16244
rect 26283 16204 26424 16232
rect 26283 16201 26295 16204
rect 26237 16195 26295 16201
rect 26418 16192 26424 16204
rect 26476 16192 26482 16244
rect 27890 16232 27896 16244
rect 27632 16204 27896 16232
rect 24026 16124 24032 16176
rect 24084 16124 24090 16176
rect 24486 16124 24492 16176
rect 24544 16124 24550 16176
rect 24688 16164 24716 16192
rect 27430 16164 27436 16176
rect 24688 16136 27436 16164
rect 22370 16096 22376 16108
rect 22066 16068 22376 16096
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 25096 16068 25237 16096
rect 25096 16056 25102 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25406 16056 25412 16108
rect 25464 16056 25470 16108
rect 26160 16105 26188 16136
rect 27430 16124 27436 16136
rect 27488 16124 27494 16176
rect 26145 16099 26203 16105
rect 26145 16065 26157 16099
rect 26191 16096 26203 16099
rect 26234 16096 26240 16108
rect 26191 16068 26240 16096
rect 26191 16065 26203 16068
rect 26145 16059 26203 16065
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 27157 16099 27215 16105
rect 27157 16065 27169 16099
rect 27203 16096 27215 16099
rect 27632 16096 27660 16204
rect 27890 16192 27896 16204
rect 27948 16232 27954 16244
rect 29365 16235 29423 16241
rect 29365 16232 29377 16235
rect 27948 16204 29377 16232
rect 27948 16192 27954 16204
rect 29365 16201 29377 16204
rect 29411 16201 29423 16235
rect 29365 16195 29423 16201
rect 28902 16124 28908 16176
rect 28960 16124 28966 16176
rect 27203 16068 27660 16096
rect 27203 16065 27215 16068
rect 27157 16059 27215 16065
rect 21174 15988 21180 16040
rect 21232 16028 21238 16040
rect 22002 16028 22008 16040
rect 21232 16000 22008 16028
rect 21232 15988 21238 16000
rect 22002 15988 22008 16000
rect 22060 16028 22066 16040
rect 22097 16031 22155 16037
rect 22097 16028 22109 16031
rect 22060 16000 22109 16028
rect 22060 15988 22066 16000
rect 22097 15997 22109 16000
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 24765 16031 24823 16037
rect 24765 15997 24777 16031
rect 24811 16028 24823 16031
rect 25130 16028 25136 16040
rect 24811 16000 25136 16028
rect 24811 15997 24823 16000
rect 24765 15991 24823 15997
rect 25130 15988 25136 16000
rect 25188 15988 25194 16040
rect 27246 15988 27252 16040
rect 27304 15988 27310 16040
rect 27614 15988 27620 16040
rect 27672 15988 27678 16040
rect 27893 16031 27951 16037
rect 27893 16028 27905 16031
rect 27724 16000 27905 16028
rect 20254 15960 20260 15972
rect 19352 15932 20260 15960
rect 20254 15920 20260 15932
rect 20312 15920 20318 15972
rect 21821 15963 21879 15969
rect 21821 15929 21833 15963
rect 21867 15960 21879 15963
rect 21910 15960 21916 15972
rect 21867 15932 21916 15960
rect 21867 15929 21879 15932
rect 21821 15923 21879 15929
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 27525 15963 27583 15969
rect 27525 15929 27537 15963
rect 27571 15960 27583 15963
rect 27724 15960 27752 16000
rect 27893 15997 27905 16000
rect 27939 15997 27951 16031
rect 27893 15991 27951 15997
rect 27571 15932 27752 15960
rect 27571 15929 27583 15932
rect 27525 15923 27583 15929
rect 9916 15864 10272 15892
rect 9916 15852 9922 15864
rect 11790 15852 11796 15904
rect 11848 15852 11854 15904
rect 12345 15895 12403 15901
rect 12345 15861 12357 15895
rect 12391 15892 12403 15895
rect 15654 15892 15660 15904
rect 12391 15864 15660 15892
rect 12391 15861 12403 15864
rect 12345 15855 12403 15861
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 17589 15895 17647 15901
rect 17589 15892 17601 15895
rect 16448 15864 17601 15892
rect 16448 15852 16454 15864
rect 17589 15861 17601 15864
rect 17635 15892 17647 15895
rect 19426 15892 19432 15904
rect 17635 15864 19432 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 19705 15895 19763 15901
rect 19705 15892 19717 15895
rect 19668 15864 19717 15892
rect 19668 15852 19674 15864
rect 19705 15861 19717 15864
rect 19751 15861 19763 15895
rect 19705 15855 19763 15861
rect 22094 15852 22100 15904
rect 22152 15852 22158 15904
rect 1104 15802 29716 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 29716 15802
rect 1104 15728 29716 15750
rect 1578 15648 1584 15700
rect 1636 15648 1642 15700
rect 2590 15648 2596 15700
rect 2648 15648 2654 15700
rect 3602 15648 3608 15700
rect 3660 15648 3666 15700
rect 3694 15648 3700 15700
rect 3752 15688 3758 15700
rect 3881 15691 3939 15697
rect 3881 15688 3893 15691
rect 3752 15660 3893 15688
rect 3752 15648 3758 15660
rect 3881 15657 3893 15660
rect 3927 15688 3939 15691
rect 4062 15688 4068 15700
rect 3927 15660 4068 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4356 15660 5304 15688
rect 4356 15620 4384 15660
rect 3436 15592 4384 15620
rect 4433 15623 4491 15629
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 2866 15484 2872 15496
rect 2556 15456 2872 15484
rect 2556 15444 2562 15456
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3326 15444 3332 15496
rect 3384 15484 3390 15496
rect 3436 15493 3464 15592
rect 4433 15589 4445 15623
rect 4479 15620 4491 15623
rect 4801 15623 4859 15629
rect 4801 15620 4813 15623
rect 4479 15592 4813 15620
rect 4479 15589 4491 15592
rect 4433 15583 4491 15589
rect 4801 15589 4813 15592
rect 4847 15589 4859 15623
rect 4801 15583 4859 15589
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 3620 15524 4721 15552
rect 3620 15493 3648 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 3421 15487 3479 15493
rect 3421 15484 3433 15487
rect 3384 15456 3433 15484
rect 3384 15444 3390 15456
rect 3421 15453 3433 15456
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3786 15444 3792 15496
rect 3844 15444 3850 15496
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 4062 15444 4068 15496
rect 4120 15484 4126 15496
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 4120 15456 4353 15484
rect 4120 15444 4126 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4614 15484 4620 15496
rect 4571 15456 4620 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4816 15484 4844 15583
rect 5166 15512 5172 15564
rect 5224 15512 5230 15564
rect 5276 15552 5304 15660
rect 5442 15648 5448 15700
rect 5500 15648 5506 15700
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 6638 15688 6644 15700
rect 6595 15660 6644 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 8938 15648 8944 15700
rect 8996 15688 9002 15700
rect 9033 15691 9091 15697
rect 9033 15688 9045 15691
rect 8996 15660 9045 15688
rect 8996 15648 9002 15660
rect 9033 15657 9045 15660
rect 9079 15657 9091 15691
rect 9033 15651 9091 15657
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10318 15688 10324 15700
rect 10100 15660 10324 15688
rect 10100 15648 10106 15660
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 10502 15648 10508 15700
rect 10560 15648 10566 15700
rect 10962 15648 10968 15700
rect 11020 15688 11026 15700
rect 11425 15691 11483 15697
rect 11425 15688 11437 15691
rect 11020 15660 11437 15688
rect 11020 15648 11026 15660
rect 11425 15657 11437 15660
rect 11471 15657 11483 15691
rect 11425 15651 11483 15657
rect 11790 15648 11796 15700
rect 11848 15648 11854 15700
rect 13262 15648 13268 15700
rect 13320 15648 13326 15700
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 16669 15691 16727 15697
rect 16669 15688 16681 15691
rect 16540 15660 16681 15688
rect 16540 15648 16546 15660
rect 16669 15657 16681 15660
rect 16715 15657 16727 15691
rect 16669 15651 16727 15657
rect 18230 15648 18236 15700
rect 18288 15688 18294 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18288 15660 18521 15688
rect 18288 15648 18294 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 18509 15651 18567 15657
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 12124 15592 13645 15620
rect 12124 15580 12130 15592
rect 13633 15589 13645 15592
rect 13679 15589 13691 15623
rect 13633 15583 13691 15589
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 5276 15524 7113 15552
rect 7101 15521 7113 15524
rect 7147 15552 7159 15555
rect 7650 15552 7656 15564
rect 7147 15524 7656 15552
rect 7147 15521 7159 15524
rect 7101 15515 7159 15521
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 9824 15524 11529 15552
rect 9824 15512 9830 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 13998 15552 14004 15564
rect 12952 15524 14004 15552
rect 12952 15512 12958 15524
rect 5184 15484 5212 15512
rect 5261 15487 5319 15493
rect 5261 15484 5273 15487
rect 4816 15456 5273 15484
rect 5261 15453 5273 15456
rect 5307 15453 5319 15487
rect 5261 15447 5319 15453
rect 5354 15487 5412 15493
rect 5354 15453 5366 15487
rect 5400 15484 5412 15487
rect 6917 15487 6975 15493
rect 5400 15456 5433 15484
rect 5400 15453 5412 15456
rect 5354 15447 5412 15453
rect 6917 15453 6929 15487
rect 6963 15484 6975 15487
rect 8478 15484 8484 15496
rect 6963 15456 8484 15484
rect 6963 15453 6975 15456
rect 6917 15447 6975 15453
rect 1486 15376 1492 15428
rect 1544 15376 1550 15428
rect 5169 15419 5227 15425
rect 5169 15385 5181 15419
rect 5215 15416 5227 15419
rect 5368 15416 5396 15447
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15484 8999 15487
rect 9030 15484 9036 15496
rect 8987 15456 9036 15484
rect 8987 15453 8999 15456
rect 8941 15447 8999 15453
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9122 15444 9128 15496
rect 9180 15444 9186 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10226 15484 10232 15496
rect 10091 15456 10232 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10226 15444 10232 15456
rect 10284 15444 10290 15496
rect 10318 15444 10324 15496
rect 10376 15444 10382 15496
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11388 15456 11437 15484
rect 11388 15444 11394 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 12986 15444 12992 15496
rect 13044 15444 13050 15496
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13170 15484 13176 15496
rect 13127 15456 13176 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13170 15444 13176 15456
rect 13228 15444 13234 15496
rect 13464 15493 13492 15524
rect 13998 15512 14004 15524
rect 14056 15552 14062 15564
rect 15286 15552 15292 15564
rect 14056 15524 14780 15552
rect 14056 15512 14062 15524
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 13541 15487 13599 15493
rect 13541 15453 13553 15487
rect 13587 15453 13599 15487
rect 13541 15447 13599 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13955 15456 14289 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 14277 15453 14289 15456
rect 14323 15484 14335 15487
rect 14366 15484 14372 15496
rect 14323 15456 14372 15484
rect 14323 15453 14335 15456
rect 14277 15447 14335 15453
rect 5626 15416 5632 15428
rect 5215 15388 5632 15416
rect 5215 15385 5227 15388
rect 5169 15379 5227 15385
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 7009 15419 7067 15425
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 7282 15416 7288 15428
rect 7055 15388 7288 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 9858 15376 9864 15428
rect 9916 15416 9922 15428
rect 10137 15419 10195 15425
rect 10137 15416 10149 15419
rect 9916 15388 10149 15416
rect 9916 15376 9922 15388
rect 10137 15385 10149 15388
rect 10183 15385 10195 15419
rect 13556 15416 13584 15447
rect 10137 15379 10195 15385
rect 10244 15388 13584 15416
rect 13740 15416 13768 15447
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14752 15416 14780 15524
rect 15028 15524 15292 15552
rect 15028 15493 15056 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 17770 15552 17776 15564
rect 15712 15524 17776 15552
rect 15712 15512 15718 15524
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 17954 15512 17960 15564
rect 18012 15512 18018 15564
rect 18524 15552 18552 15651
rect 18874 15648 18880 15700
rect 18932 15688 18938 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 18932 15660 19717 15688
rect 18932 15648 18938 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 19981 15691 20039 15697
rect 19981 15657 19993 15691
rect 20027 15688 20039 15691
rect 20346 15688 20352 15700
rect 20027 15660 20352 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 21266 15688 21272 15700
rect 21039 15660 21272 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 22278 15620 22284 15632
rect 22112 15592 22284 15620
rect 19337 15555 19395 15561
rect 19337 15552 19349 15555
rect 18524 15524 19349 15552
rect 19337 15521 19349 15524
rect 19383 15521 19395 15555
rect 19337 15515 19395 15521
rect 19886 15512 19892 15564
rect 19944 15552 19950 15564
rect 22112 15561 22140 15592
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 20809 15555 20867 15561
rect 20809 15552 20821 15555
rect 19944 15524 20821 15552
rect 19944 15512 19950 15524
rect 20809 15521 20821 15524
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 22097 15555 22155 15561
rect 22097 15521 22109 15555
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 23753 15555 23811 15561
rect 23753 15552 23765 15555
rect 23624 15524 23765 15552
rect 23624 15512 23630 15524
rect 23753 15521 23765 15524
rect 23799 15521 23811 15555
rect 23753 15515 23811 15521
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15484 15255 15487
rect 16298 15484 16304 15496
rect 15243 15456 16304 15484
rect 15243 15453 15255 15456
rect 15197 15447 15255 15453
rect 15212 15416 15240 15447
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 17310 15444 17316 15496
rect 17368 15444 17374 15496
rect 17494 15444 17500 15496
rect 17552 15444 17558 15496
rect 17586 15444 17592 15496
rect 17644 15444 17650 15496
rect 17681 15487 17739 15493
rect 17681 15453 17693 15487
rect 17727 15484 17739 15487
rect 17788 15484 17816 15512
rect 17727 15456 17816 15484
rect 18049 15487 18107 15493
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 18049 15453 18061 15487
rect 18095 15453 18107 15487
rect 18049 15447 18107 15453
rect 18141 15487 18199 15493
rect 18141 15453 18153 15487
rect 18187 15484 18199 15487
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18187 15456 18337 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 13740 15388 14504 15416
rect 14752 15388 15240 15416
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 10244 15348 10272 15388
rect 9824 15320 10272 15348
rect 9824 15308 9830 15320
rect 12618 15308 12624 15360
rect 12676 15308 12682 15360
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 14274 15348 14280 15360
rect 13136 15320 14280 15348
rect 13136 15308 13142 15320
rect 14274 15308 14280 15320
rect 14332 15348 14338 15360
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 14332 15320 14381 15348
rect 14332 15308 14338 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14476 15348 14504 15388
rect 15286 15376 15292 15428
rect 15344 15416 15350 15428
rect 15381 15419 15439 15425
rect 15381 15416 15393 15419
rect 15344 15388 15393 15416
rect 15344 15376 15350 15388
rect 15381 15385 15393 15388
rect 15427 15385 15439 15419
rect 17328 15416 17356 15444
rect 18064 15416 18092 15447
rect 17328 15388 18092 15416
rect 15381 15379 15439 15385
rect 18230 15376 18236 15428
rect 18288 15416 18294 15428
rect 18524 15416 18552 15447
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19797 15487 19855 15493
rect 19797 15484 19809 15487
rect 19576 15456 19809 15484
rect 19576 15444 19582 15456
rect 19797 15453 19809 15456
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 20714 15444 20720 15496
rect 20772 15444 20778 15496
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 22189 15487 22247 15493
rect 22189 15453 22201 15487
rect 22235 15484 22247 15487
rect 22370 15484 22376 15496
rect 22235 15456 22376 15484
rect 22235 15453 22247 15456
rect 22189 15447 22247 15453
rect 18288 15388 18552 15416
rect 21008 15416 21036 15447
rect 22370 15444 22376 15456
rect 22428 15444 22434 15496
rect 23658 15484 23664 15496
rect 22480 15456 23664 15484
rect 21008 15388 21957 15416
rect 18288 15376 18294 15388
rect 21177 15351 21235 15357
rect 21177 15348 21189 15351
rect 14476 15320 21189 15348
rect 14369 15311 14427 15317
rect 21177 15317 21189 15320
rect 21223 15317 21235 15351
rect 21929 15348 21957 15388
rect 22002 15376 22008 15428
rect 22060 15416 22066 15428
rect 22480 15416 22508 15456
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15484 24639 15487
rect 24670 15484 24676 15496
rect 24627 15456 24676 15484
rect 24627 15453 24639 15456
rect 24581 15447 24639 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 27338 15444 27344 15496
rect 27396 15444 27402 15496
rect 27525 15487 27583 15493
rect 27525 15453 27537 15487
rect 27571 15453 27583 15487
rect 27525 15447 27583 15453
rect 23569 15419 23627 15425
rect 23569 15416 23581 15419
rect 22060 15388 22508 15416
rect 22572 15388 23581 15416
rect 22060 15376 22066 15388
rect 22462 15348 22468 15360
rect 21929 15320 22468 15348
rect 21177 15311 21235 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 22572 15357 22600 15388
rect 23569 15385 23581 15388
rect 23615 15385 23627 15419
rect 23569 15379 23627 15385
rect 27154 15376 27160 15428
rect 27212 15416 27218 15428
rect 27540 15416 27568 15447
rect 29086 15444 29092 15496
rect 29144 15444 29150 15496
rect 29362 15444 29368 15496
rect 29420 15444 29426 15496
rect 27212 15388 27568 15416
rect 27212 15376 27218 15388
rect 22557 15351 22615 15357
rect 22557 15317 22569 15351
rect 22603 15317 22615 15351
rect 22557 15311 22615 15317
rect 23198 15308 23204 15360
rect 23256 15308 23262 15360
rect 24394 15308 24400 15360
rect 24452 15348 24458 15360
rect 24489 15351 24547 15357
rect 24489 15348 24501 15351
rect 24452 15320 24501 15348
rect 24452 15308 24458 15320
rect 24489 15317 24501 15320
rect 24535 15317 24547 15351
rect 24489 15311 24547 15317
rect 27246 15308 27252 15360
rect 27304 15348 27310 15360
rect 27433 15351 27491 15357
rect 27433 15348 27445 15351
rect 27304 15320 27445 15348
rect 27304 15308 27310 15320
rect 27433 15317 27445 15320
rect 27479 15348 27491 15351
rect 28534 15348 28540 15360
rect 27479 15320 28540 15348
rect 27479 15317 27491 15320
rect 27433 15311 27491 15317
rect 28534 15308 28540 15320
rect 28592 15308 28598 15360
rect 1104 15258 29716 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 29716 15258
rect 1104 15184 29716 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 9674 15144 9680 15156
rect 4120 15116 9680 15144
rect 4120 15104 4126 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 11606 15144 11612 15156
rect 10192 15116 11612 15144
rect 10192 15104 10198 15116
rect 11606 15104 11612 15116
rect 11664 15144 11670 15156
rect 12342 15144 12348 15156
rect 11664 15116 12348 15144
rect 11664 15104 11670 15116
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12713 15147 12771 15153
rect 12713 15144 12725 15147
rect 12676 15116 12725 15144
rect 12676 15104 12682 15116
rect 12713 15113 12725 15116
rect 12759 15113 12771 15147
rect 12713 15107 12771 15113
rect 12986 15104 12992 15156
rect 13044 15144 13050 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 13044 15116 13369 15144
rect 13044 15104 13050 15116
rect 13357 15113 13369 15116
rect 13403 15113 13415 15147
rect 13357 15107 13415 15113
rect 16945 15147 17003 15153
rect 16945 15113 16957 15147
rect 16991 15144 17003 15147
rect 17310 15144 17316 15156
rect 16991 15116 17316 15144
rect 16991 15113 17003 15116
rect 16945 15107 17003 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 20898 15144 20904 15156
rect 19300 15116 20904 15144
rect 19300 15104 19306 15116
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 27890 15144 27896 15156
rect 23716 15116 25084 15144
rect 23716 15104 23722 15116
rect 6656 15048 6960 15076
rect 6656 15020 6684 15048
rect 6638 14968 6644 15020
rect 6696 14968 6702 15020
rect 6932 15017 6960 15048
rect 7834 15036 7840 15088
rect 7892 15076 7898 15088
rect 16206 15076 16212 15088
rect 7892 15048 13400 15076
rect 15778 15048 16212 15076
rect 7892 15036 7898 15048
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 6917 14971 6975 14977
rect 6840 14940 6868 14971
rect 7098 14968 7104 15020
rect 7156 14968 7162 15020
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 11146 14968 11152 15020
rect 11204 15008 11210 15020
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 11204 14980 11529 15008
rect 11204 14968 11210 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 11517 14971 11575 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 11992 15017 12020 15048
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11664 14980 11713 15008
rect 11664 14968 11670 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 12342 14968 12348 15020
rect 12400 14968 12406 15020
rect 12434 14968 12440 15020
rect 12492 14968 12498 15020
rect 13004 15017 13032 15048
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 7116 14940 7144 14968
rect 6840 14912 7144 14940
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 12912 14940 12940 14971
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 13372 15017 13400 15048
rect 16206 15036 16212 15048
rect 16264 15036 16270 15088
rect 16298 15036 16304 15088
rect 16356 15036 16362 15088
rect 19334 15076 19340 15088
rect 17052 15048 19340 15076
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 14977 13599 15011
rect 16316 15008 16344 15036
rect 17052 15017 17080 15048
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 23198 15036 23204 15088
rect 23256 15076 23262 15088
rect 25056 15085 25084 15116
rect 27264 15116 27896 15144
rect 23293 15079 23351 15085
rect 23293 15076 23305 15079
rect 23256 15048 23305 15076
rect 23256 15036 23262 15048
rect 23293 15045 23305 15048
rect 23339 15045 23351 15079
rect 23293 15039 23351 15045
rect 25041 15079 25099 15085
rect 25041 15045 25053 15079
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 16316 14980 16773 15008
rect 13541 14971 13599 14977
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 15008 17003 15011
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16991 14980 17049 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17037 14971 17095 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17402 15008 17408 15020
rect 17267 14980 17408 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 13078 14940 13084 14952
rect 8352 14912 12020 14940
rect 12912 14912 13084 14940
rect 8352 14900 8358 14912
rect 1946 14832 1952 14884
rect 2004 14872 2010 14884
rect 9122 14872 9128 14884
rect 2004 14844 9128 14872
rect 2004 14832 2010 14844
rect 9122 14832 9128 14844
rect 9180 14832 9186 14884
rect 11882 14832 11888 14884
rect 11940 14832 11946 14884
rect 11992 14872 12020 14912
rect 13078 14900 13084 14912
rect 13136 14940 13142 14952
rect 13556 14940 13584 14971
rect 13136 14912 13584 14940
rect 13136 14900 13142 14912
rect 14274 14900 14280 14952
rect 14332 14900 14338 14952
rect 14550 14900 14556 14952
rect 14608 14900 14614 14952
rect 16776 14940 16804 14971
rect 17236 14940 17264 14971
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 22002 14968 22008 15020
rect 22060 14968 22066 15020
rect 24394 14968 24400 15020
rect 24452 14968 24458 15020
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 15008 26203 15011
rect 26234 15008 26240 15020
rect 26191 14980 26240 15008
rect 26191 14977 26203 14980
rect 26145 14971 26203 14977
rect 26234 14968 26240 14980
rect 26292 14968 26298 15020
rect 27264 15017 27292 15116
rect 27890 15104 27896 15116
rect 27948 15104 27954 15156
rect 27982 15104 27988 15156
rect 28040 15144 28046 15156
rect 28040 15116 28488 15144
rect 28040 15104 28046 15116
rect 27801 15079 27859 15085
rect 27801 15045 27813 15079
rect 27847 15076 27859 15079
rect 27847 15048 28120 15076
rect 27847 15045 27859 15048
rect 27801 15039 27859 15045
rect 27249 15011 27307 15017
rect 27249 14977 27261 15011
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 27985 15011 28043 15017
rect 27985 14977 27997 15011
rect 28031 14977 28043 15011
rect 27985 14971 28043 14977
rect 16776 14912 17264 14940
rect 20898 14900 20904 14952
rect 20956 14940 20962 14952
rect 21913 14943 21971 14949
rect 21913 14940 21925 14943
rect 20956 14912 21925 14940
rect 20956 14900 20962 14912
rect 21913 14909 21925 14912
rect 21959 14909 21971 14943
rect 21913 14903 21971 14909
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 22336 14912 22385 14940
rect 22336 14900 22342 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 23017 14943 23075 14949
rect 23017 14909 23029 14943
rect 23063 14940 23075 14943
rect 25130 14940 25136 14952
rect 23063 14912 25136 14940
rect 23063 14909 23075 14912
rect 23017 14903 23075 14909
rect 25130 14900 25136 14912
rect 25188 14900 25194 14952
rect 25869 14943 25927 14949
rect 25869 14909 25881 14943
rect 25915 14940 25927 14943
rect 26050 14940 26056 14952
rect 25915 14912 26056 14940
rect 25915 14909 25927 14912
rect 25869 14903 25927 14909
rect 26050 14900 26056 14912
rect 26108 14940 26114 14952
rect 26108 14912 27108 14940
rect 26108 14900 26114 14912
rect 12434 14872 12440 14884
rect 11992 14844 12440 14872
rect 12434 14832 12440 14844
rect 12492 14832 12498 14884
rect 13173 14875 13231 14881
rect 13173 14841 13185 14875
rect 13219 14872 13231 14875
rect 13538 14872 13544 14884
rect 13219 14844 13544 14872
rect 13219 14841 13231 14844
rect 13173 14835 13231 14841
rect 13538 14832 13544 14844
rect 13596 14872 13602 14884
rect 14090 14872 14096 14884
rect 13596 14844 14096 14872
rect 13596 14832 13602 14844
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 22922 14872 22928 14884
rect 15580 14844 22928 14872
rect 6730 14764 6736 14816
rect 6788 14764 6794 14816
rect 6914 14764 6920 14816
rect 6972 14764 6978 14816
rect 10045 14807 10103 14813
rect 10045 14773 10057 14807
rect 10091 14804 10103 14807
rect 10134 14804 10140 14816
rect 10091 14776 10140 14804
rect 10091 14773 10103 14776
rect 10045 14767 10103 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 12452 14804 12480 14832
rect 13262 14804 13268 14816
rect 12452 14776 13268 14804
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 15580 14804 15608 14844
rect 22922 14832 22928 14844
rect 22980 14832 22986 14884
rect 25593 14875 25651 14881
rect 25593 14841 25605 14875
rect 25639 14872 25651 14875
rect 26973 14875 27031 14881
rect 26973 14872 26985 14875
rect 25639 14844 26985 14872
rect 25639 14841 25651 14844
rect 25593 14835 25651 14841
rect 26973 14841 26985 14844
rect 27019 14841 27031 14875
rect 26973 14835 27031 14841
rect 13412 14776 15608 14804
rect 17221 14807 17279 14813
rect 13412 14764 13418 14776
rect 17221 14773 17233 14807
rect 17267 14804 17279 14807
rect 18230 14804 18236 14816
rect 17267 14776 18236 14804
rect 17267 14773 17279 14776
rect 17221 14767 17279 14773
rect 18230 14764 18236 14776
rect 18288 14764 18294 14816
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 22094 14804 22100 14816
rect 20496 14776 22100 14804
rect 20496 14764 20502 14776
rect 22094 14764 22100 14776
rect 22152 14764 22158 14816
rect 25406 14764 25412 14816
rect 25464 14764 25470 14816
rect 26053 14807 26111 14813
rect 26053 14773 26065 14807
rect 26099 14804 26111 14807
rect 26234 14804 26240 14816
rect 26099 14776 26240 14804
rect 26099 14773 26111 14776
rect 26053 14767 26111 14773
rect 26234 14764 26240 14776
rect 26292 14764 26298 14816
rect 27080 14804 27108 14912
rect 27154 14900 27160 14952
rect 27212 14900 27218 14952
rect 27338 14900 27344 14952
rect 27396 14900 27402 14952
rect 27430 14900 27436 14952
rect 27488 14940 27494 14952
rect 28000 14940 28028 14971
rect 27488 14912 28028 14940
rect 27488 14900 27494 14912
rect 27172 14872 27200 14900
rect 28092 14872 28120 15048
rect 28460 15017 28488 15116
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 28534 14968 28540 15020
rect 28592 14968 28598 15020
rect 27172 14844 28120 14872
rect 28166 14832 28172 14884
rect 28224 14872 28230 14884
rect 28224 14844 29776 14872
rect 28224 14832 28230 14844
rect 27617 14807 27675 14813
rect 27617 14804 27629 14807
rect 27080 14776 27629 14804
rect 27617 14773 27629 14776
rect 27663 14773 27675 14807
rect 27617 14767 27675 14773
rect 28258 14764 28264 14816
rect 28316 14764 28322 14816
rect 1104 14714 29716 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 29716 14714
rect 1104 14640 29716 14662
rect 6730 14560 6736 14612
rect 6788 14560 6794 14612
rect 6822 14560 6828 14612
rect 6880 14600 6886 14612
rect 14182 14600 14188 14612
rect 6880 14572 14188 14600
rect 6880 14560 6886 14572
rect 6365 14535 6423 14541
rect 6365 14501 6377 14535
rect 6411 14532 6423 14535
rect 6914 14532 6920 14544
rect 6411 14504 6920 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4798 14464 4804 14476
rect 4479 14436 4804 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4798 14424 4804 14436
rect 4856 14464 4862 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 4856 14436 7021 14464
rect 4856 14424 4862 14436
rect 7009 14433 7021 14436
rect 7055 14464 7067 14467
rect 7374 14464 7380 14476
rect 7055 14436 7380 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 8536 14436 8769 14464
rect 8536 14424 8542 14436
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 2774 14356 2780 14408
rect 2832 14396 2838 14408
rect 3421 14399 3479 14405
rect 3421 14396 3433 14399
rect 2832 14368 3433 14396
rect 2832 14356 2838 14368
rect 3421 14365 3433 14368
rect 3467 14365 3479 14399
rect 3421 14359 3479 14365
rect 5994 14356 6000 14408
rect 6052 14396 6058 14408
rect 6822 14396 6828 14408
rect 6052 14368 6828 14396
rect 6052 14356 6058 14368
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 9140 14405 9168 14572
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 14550 14600 14556 14612
rect 14323 14572 14556 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 14550 14560 14556 14572
rect 14608 14560 14614 14612
rect 15930 14560 15936 14612
rect 15988 14560 15994 14612
rect 16206 14560 16212 14612
rect 16264 14560 16270 14612
rect 26605 14603 26663 14609
rect 16316 14572 26188 14600
rect 10042 14492 10048 14544
rect 10100 14532 10106 14544
rect 10318 14532 10324 14544
rect 10100 14504 10324 14532
rect 10100 14492 10106 14504
rect 10318 14492 10324 14504
rect 10376 14532 10382 14544
rect 10594 14532 10600 14544
rect 10376 14504 10600 14532
rect 10376 14492 10382 14504
rect 10594 14492 10600 14504
rect 10652 14532 10658 14544
rect 10652 14504 10916 14532
rect 10652 14492 10658 14504
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 10778 14464 10784 14476
rect 9272 14436 10784 14464
rect 9272 14424 9278 14436
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 10888 14464 10916 14504
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 16316 14532 16344 14572
rect 11296 14504 16344 14532
rect 11296 14492 11302 14504
rect 17954 14492 17960 14544
rect 18012 14492 18018 14544
rect 18049 14535 18107 14541
rect 18049 14501 18061 14535
rect 18095 14532 18107 14535
rect 18230 14532 18236 14544
rect 18095 14504 18236 14532
rect 18095 14501 18107 14504
rect 18049 14495 18107 14501
rect 18230 14492 18236 14504
rect 18288 14492 18294 14544
rect 18506 14492 18512 14544
rect 18564 14532 18570 14544
rect 19337 14535 19395 14541
rect 19337 14532 19349 14535
rect 18564 14504 19349 14532
rect 18564 14492 18570 14504
rect 19337 14501 19349 14504
rect 19383 14532 19395 14535
rect 19518 14532 19524 14544
rect 19383 14504 19524 14532
rect 19383 14501 19395 14504
rect 19337 14495 19395 14501
rect 19518 14492 19524 14504
rect 19576 14492 19582 14544
rect 13449 14467 13507 14473
rect 10888 14436 13400 14464
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 10042 14356 10048 14408
rect 10100 14356 10106 14408
rect 10134 14356 10140 14408
rect 10192 14396 10198 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10192 14368 10425 14396
rect 10192 14356 10198 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10594 14356 10600 14408
rect 10652 14356 10658 14408
rect 10965 14399 11023 14405
rect 10965 14365 10977 14399
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13136 14368 13185 14396
rect 13136 14356 13142 14368
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13372 14396 13400 14436
rect 13449 14433 13461 14467
rect 13495 14464 13507 14467
rect 13998 14464 14004 14476
rect 13495 14436 14004 14464
rect 13495 14433 13507 14436
rect 13449 14427 13507 14433
rect 13998 14424 14004 14436
rect 14056 14424 14062 14476
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 15010 14464 15016 14476
rect 14240 14436 15016 14464
rect 14240 14424 14246 14436
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14464 15807 14467
rect 16390 14464 16396 14476
rect 15795 14436 16396 14464
rect 15795 14433 15807 14436
rect 15749 14427 15807 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 17972 14464 18000 14492
rect 17512 14436 18000 14464
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 13372 14368 13645 14396
rect 13265 14359 13323 14365
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 4706 14288 4712 14340
rect 4764 14288 4770 14340
rect 5442 14288 5448 14340
rect 5500 14288 5506 14340
rect 6362 14328 6368 14340
rect 6104 14300 6368 14328
rect 3418 14220 3424 14272
rect 3476 14260 3482 14272
rect 3513 14263 3571 14269
rect 3513 14260 3525 14263
rect 3476 14232 3525 14260
rect 3476 14220 3482 14232
rect 3513 14229 3525 14232
rect 3559 14229 3571 14263
rect 3513 14223 3571 14229
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 6104 14260 6132 14300
rect 6362 14288 6368 14300
rect 6420 14328 6426 14340
rect 6733 14331 6791 14337
rect 6733 14328 6745 14331
rect 6420 14300 6745 14328
rect 6420 14288 6426 14300
rect 6733 14297 6745 14300
rect 6779 14297 6791 14331
rect 7285 14331 7343 14337
rect 7285 14328 7297 14331
rect 6733 14291 6791 14297
rect 6932 14300 7297 14328
rect 5592 14232 6132 14260
rect 5592 14220 5598 14232
rect 6178 14220 6184 14272
rect 6236 14220 6242 14272
rect 6932 14269 6960 14300
rect 7285 14297 7297 14300
rect 7331 14297 7343 14331
rect 9033 14331 9091 14337
rect 9033 14328 9045 14331
rect 8510 14300 9045 14328
rect 7285 14291 7343 14297
rect 9033 14297 9045 14300
rect 9079 14297 9091 14331
rect 9033 14291 9091 14297
rect 10321 14331 10379 14337
rect 10321 14297 10333 14331
rect 10367 14328 10379 14331
rect 11514 14328 11520 14340
rect 10367 14300 11520 14328
rect 10367 14297 10379 14300
rect 10321 14291 10379 14297
rect 10612 14272 10640 14300
rect 11514 14288 11520 14300
rect 11572 14288 11578 14340
rect 12986 14288 12992 14340
rect 13044 14328 13050 14340
rect 13280 14328 13308 14359
rect 13044 14300 13308 14328
rect 13648 14328 13676 14359
rect 13814 14356 13820 14408
rect 13872 14356 13878 14408
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14461 14399 14519 14405
rect 14461 14396 14473 14399
rect 14424 14368 14473 14396
rect 14424 14356 14430 14368
rect 14461 14365 14473 14368
rect 14507 14365 14519 14399
rect 14461 14359 14519 14365
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14396 14795 14399
rect 15194 14396 15200 14408
rect 14783 14368 15200 14396
rect 14783 14365 14795 14368
rect 14737 14359 14795 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 17512 14405 17540 14436
rect 18322 14424 18328 14476
rect 18380 14424 18386 14476
rect 18598 14424 18604 14476
rect 18656 14424 18662 14476
rect 19061 14467 19119 14473
rect 19061 14433 19073 14467
rect 19107 14464 19119 14467
rect 20070 14464 20076 14476
rect 19107 14436 20076 14464
rect 19107 14433 19119 14436
rect 19061 14427 19119 14433
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 24857 14467 24915 14473
rect 24857 14433 24869 14467
rect 24903 14464 24915 14467
rect 25130 14464 25136 14476
rect 24903 14436 25136 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 25130 14424 25136 14436
rect 25188 14424 25194 14476
rect 26160 14464 26188 14572
rect 26605 14569 26617 14603
rect 26651 14600 26663 14603
rect 27430 14600 27436 14612
rect 26651 14572 27436 14600
rect 26651 14569 26663 14572
rect 26605 14563 26663 14569
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 27525 14603 27583 14609
rect 27525 14569 27537 14603
rect 27571 14600 27583 14603
rect 27706 14600 27712 14612
rect 27571 14572 27712 14600
rect 27571 14569 27583 14572
rect 27525 14563 27583 14569
rect 27706 14560 27712 14572
rect 27764 14560 27770 14612
rect 27880 14603 27938 14609
rect 27880 14569 27892 14603
rect 27926 14600 27938 14603
rect 28258 14600 28264 14612
rect 27926 14572 28264 14600
rect 27926 14569 27938 14572
rect 27880 14563 27938 14569
rect 28258 14560 28264 14572
rect 28316 14560 28322 14612
rect 29365 14603 29423 14609
rect 29365 14569 29377 14603
rect 29411 14600 29423 14603
rect 29748 14600 29776 14844
rect 29411 14572 29776 14600
rect 29411 14569 29423 14572
rect 29365 14563 29423 14569
rect 29086 14464 29092 14476
rect 26160 14436 29092 14464
rect 29086 14424 29092 14436
rect 29144 14424 29150 14476
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14365 16359 14399
rect 16301 14359 16359 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14365 17739 14399
rect 17681 14359 17739 14365
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 14550 14328 14556 14340
rect 13648 14300 14556 14328
rect 13044 14288 13050 14300
rect 14550 14288 14556 14300
rect 14608 14288 14614 14340
rect 15010 14288 15016 14340
rect 15068 14328 15074 14340
rect 16316 14328 16344 14359
rect 17034 14328 17040 14340
rect 15068 14300 17040 14328
rect 15068 14288 15074 14300
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14229 6975 14263
rect 6917 14223 6975 14229
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10870 14220 10876 14272
rect 10928 14220 10934 14272
rect 13446 14220 13452 14272
rect 13504 14220 13510 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 13725 14263 13783 14269
rect 13725 14260 13737 14263
rect 13688 14232 13737 14260
rect 13688 14220 13694 14232
rect 13725 14229 13737 14232
rect 13771 14229 13783 14263
rect 13725 14223 13783 14229
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17589 14263 17647 14269
rect 17589 14260 17601 14263
rect 17460 14232 17601 14260
rect 17460 14220 17466 14232
rect 17589 14229 17601 14232
rect 17635 14229 17647 14263
rect 17696 14260 17724 14359
rect 17880 14328 17908 14359
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18506 14396 18512 14408
rect 18196 14368 18512 14396
rect 18196 14356 18202 14368
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 18874 14396 18880 14408
rect 18739 14368 18880 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18874 14356 18880 14368
rect 18932 14356 18938 14408
rect 19245 14399 19303 14405
rect 19245 14365 19257 14399
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 18322 14328 18328 14340
rect 17880 14300 18328 14328
rect 18322 14288 18328 14300
rect 18380 14328 18386 14340
rect 19260 14328 19288 14359
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 19702 14356 19708 14408
rect 19760 14356 19766 14408
rect 26234 14356 26240 14408
rect 26292 14356 26298 14408
rect 27614 14356 27620 14408
rect 27672 14356 27678 14408
rect 18380 14300 19288 14328
rect 18380 14288 18386 14300
rect 19978 14288 19984 14340
rect 20036 14288 20042 14340
rect 20990 14288 20996 14340
rect 21048 14288 21054 14340
rect 21729 14331 21787 14337
rect 21729 14297 21741 14331
rect 21775 14297 21787 14331
rect 21729 14291 21787 14297
rect 25133 14331 25191 14337
rect 25133 14297 25145 14331
rect 25179 14328 25191 14331
rect 25406 14328 25412 14340
rect 25179 14300 25412 14328
rect 25179 14297 25191 14300
rect 25133 14291 25191 14297
rect 18230 14260 18236 14272
rect 17696 14232 18236 14260
rect 17589 14223 17647 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 20254 14220 20260 14272
rect 20312 14260 20318 14272
rect 21744 14260 21772 14291
rect 25406 14288 25412 14300
rect 25464 14288 25470 14340
rect 27154 14288 27160 14340
rect 27212 14288 27218 14340
rect 27338 14288 27344 14340
rect 27396 14328 27402 14340
rect 28166 14328 28172 14340
rect 27396 14300 28172 14328
rect 27396 14288 27402 14300
rect 28166 14288 28172 14300
rect 28224 14288 28230 14340
rect 28902 14288 28908 14340
rect 28960 14288 28966 14340
rect 20312 14232 21772 14260
rect 20312 14220 20318 14232
rect 22278 14220 22284 14272
rect 22336 14260 22342 14272
rect 29178 14260 29184 14272
rect 22336 14232 29184 14260
rect 22336 14220 22342 14232
rect 29178 14220 29184 14232
rect 29236 14220 29242 14272
rect 1104 14170 29716 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 29716 14170
rect 1104 14096 29716 14118
rect 4798 14056 4804 14068
rect 2424 14028 4804 14056
rect 1394 13812 1400 13864
rect 1452 13812 1458 13864
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 1719 13824 1900 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1872 13784 1900 13824
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 2424 13861 2452 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5442 14016 5448 14068
rect 5500 14016 5506 14068
rect 6178 14016 6184 14068
rect 6236 14056 6242 14068
rect 7006 14056 7012 14068
rect 6236 14028 7012 14056
rect 6236 14016 6242 14028
rect 3418 13948 3424 14000
rect 3476 13948 3482 14000
rect 4709 13991 4767 13997
rect 4709 13957 4721 13991
rect 4755 13988 4767 13991
rect 5534 13988 5540 14000
rect 4755 13960 5540 13988
rect 4755 13957 4767 13960
rect 4709 13951 4767 13957
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 6564 13997 6592 14028
rect 7006 14016 7012 14028
rect 7064 14056 7070 14068
rect 10318 14056 10324 14068
rect 7064 14028 10324 14056
rect 7064 14016 7070 14028
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 12158 14016 12164 14068
rect 12216 14016 12222 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14025 12311 14059
rect 16025 14059 16083 14065
rect 12253 14019 12311 14025
rect 13740 14028 14688 14056
rect 6549 13991 6607 13997
rect 6549 13957 6561 13991
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 6914 13988 6920 14000
rect 6779 13960 6920 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 9401 13991 9459 13997
rect 9401 13988 9413 13991
rect 9140 13960 9413 13988
rect 9140 13932 9168 13960
rect 9401 13957 9413 13960
rect 9447 13957 9459 13991
rect 9401 13951 9459 13957
rect 9493 13991 9551 13997
rect 9493 13957 9505 13991
rect 9539 13988 9551 13991
rect 10873 13991 10931 13997
rect 9539 13960 10456 13988
rect 9539 13957 9551 13960
rect 9493 13951 9551 13957
rect 4614 13880 4620 13932
rect 4672 13920 4678 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4672 13892 5089 13920
rect 4672 13880 4678 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 5353 13923 5411 13929
rect 5353 13889 5365 13923
rect 5399 13920 5411 13923
rect 5442 13920 5448 13932
rect 5399 13892 5448 13920
rect 5399 13889 5411 13892
rect 5353 13883 5411 13889
rect 5442 13880 5448 13892
rect 5500 13920 5506 13932
rect 5994 13920 6000 13932
rect 5500 13892 6000 13920
rect 5500 13880 5506 13892
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6822 13880 6828 13932
rect 6880 13880 6886 13932
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 7392 13892 7481 13920
rect 2409 13855 2467 13861
rect 2409 13852 2421 13855
rect 2004 13824 2421 13852
rect 2004 13812 2010 13824
rect 2409 13821 2421 13824
rect 2455 13821 2467 13855
rect 4062 13852 4068 13864
rect 2409 13815 2467 13821
rect 2516 13824 4068 13852
rect 2516 13784 2544 13824
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4706 13852 4712 13864
rect 4540 13824 4712 13852
rect 4540 13793 4568 13824
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 7190 13812 7196 13864
rect 7248 13852 7254 13864
rect 7392 13852 7420 13892
rect 7469 13889 7481 13892
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 8294 13920 8300 13932
rect 7607 13892 8300 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 9122 13880 9128 13932
rect 9180 13880 9186 13932
rect 9214 13880 9220 13932
rect 9272 13880 9278 13932
rect 9508 13852 9536 13951
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 7248 13824 7420 13852
rect 8036 13824 9536 13852
rect 7248 13812 7254 13824
rect 1872 13756 2544 13784
rect 4525 13787 4583 13793
rect 4525 13753 4537 13787
rect 4571 13753 4583 13787
rect 6365 13787 6423 13793
rect 6365 13784 6377 13787
rect 4525 13747 4583 13753
rect 5368 13756 6377 13784
rect 2672 13719 2730 13725
rect 2672 13685 2684 13719
rect 2718 13716 2730 13719
rect 3786 13716 3792 13728
rect 2718 13688 3792 13716
rect 2718 13685 2730 13688
rect 2672 13679 2730 13685
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 4120 13688 4169 13716
rect 4120 13676 4126 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4157 13679 4215 13685
rect 4709 13719 4767 13725
rect 4709 13685 4721 13719
rect 4755 13716 4767 13719
rect 5368 13716 5396 13756
rect 6365 13753 6377 13756
rect 6411 13753 6423 13787
rect 6365 13747 6423 13753
rect 4755 13688 5396 13716
rect 6917 13719 6975 13725
rect 4755 13685 4767 13688
rect 4709 13679 4767 13685
rect 6917 13685 6929 13719
rect 6963 13716 6975 13719
rect 7098 13716 7104 13728
rect 6963 13688 7104 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 7098 13676 7104 13688
rect 7156 13716 7162 13728
rect 8036 13716 8064 13824
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 9600 13784 9628 13883
rect 10428 13852 10456 13960
rect 10873 13957 10885 13991
rect 10919 13988 10931 13991
rect 11238 13988 11244 14000
rect 10919 13960 11244 13988
rect 10919 13957 10931 13960
rect 10873 13951 10931 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 11606 13988 11612 14000
rect 11440 13960 11612 13988
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10778 13929 10784 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10560 13892 10609 13920
rect 10560 13880 10566 13892
rect 10597 13889 10609 13892
rect 10643 13889 10655 13923
rect 10597 13883 10655 13889
rect 10745 13923 10784 13929
rect 10745 13889 10757 13923
rect 10745 13883 10784 13889
rect 10612 13852 10640 13883
rect 10778 13880 10784 13883
rect 10836 13880 10842 13932
rect 10962 13880 10968 13932
rect 11020 13880 11026 13932
rect 11054 13880 11060 13932
rect 11112 13929 11118 13932
rect 11112 13923 11161 13929
rect 11112 13889 11115 13923
rect 11149 13920 11161 13923
rect 11440 13920 11468 13960
rect 11606 13948 11612 13960
rect 11664 13948 11670 14000
rect 12002 13991 12060 13997
rect 12002 13957 12014 13991
rect 12048 13988 12060 13991
rect 12268 13988 12296 14019
rect 12048 13960 12296 13988
rect 12048 13957 12060 13960
rect 12002 13951 12060 13957
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13740 13988 13768 14028
rect 13136 13960 13768 13988
rect 13136 13948 13142 13960
rect 11149 13892 11468 13920
rect 11149 13889 11161 13892
rect 11112 13883 11161 13889
rect 11112 13880 11118 13883
rect 11514 13880 11520 13932
rect 11572 13880 11578 13932
rect 12986 13929 12992 13932
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 11624 13892 12633 13920
rect 11624 13852 11652 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12943 13923 12992 13929
rect 12943 13920 12955 13923
rect 12621 13883 12679 13889
rect 12728 13892 12955 13920
rect 10428 13824 10548 13852
rect 10612 13824 11652 13852
rect 10410 13784 10416 13796
rect 8260 13756 10416 13784
rect 8260 13744 8266 13756
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 10520 13784 10548 13824
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12434 13852 12440 13864
rect 11931 13824 12440 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 12728 13852 12756 13892
rect 12943 13889 12955 13892
rect 12989 13889 12992 13923
rect 12943 13883 12992 13889
rect 12986 13880 12992 13883
rect 13044 13880 13050 13932
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13354 13920 13360 13932
rect 13315 13892 13360 13920
rect 13173 13883 13231 13889
rect 12575 13824 12756 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 10962 13784 10968 13796
rect 10520 13756 10968 13784
rect 10962 13744 10968 13756
rect 11020 13784 11026 13796
rect 12544 13784 12572 13815
rect 11020 13756 12572 13784
rect 13004 13784 13032 13880
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 13188 13852 13216 13883
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 13630 13920 13636 13932
rect 13495 13892 13636 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13740 13929 13768 13960
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 14277 13991 14335 13997
rect 14277 13988 14289 13991
rect 13872 13960 14289 13988
rect 13872 13948 13878 13960
rect 14277 13957 14289 13960
rect 14323 13988 14335 13991
rect 14323 13960 14504 13988
rect 14323 13957 14335 13960
rect 14277 13951 14335 13957
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 13998 13880 14004 13932
rect 14056 13880 14062 13932
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14476 13929 14504 13960
rect 14550 13948 14556 14000
rect 14608 13948 14614 14000
rect 14660 13988 14688 14028
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 16071 14028 16957 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 16945 14019 17003 14025
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18877 14059 18935 14065
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 19426 14056 19432 14068
rect 18923 14028 19432 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 19978 14056 19984 14068
rect 19843 14028 19984 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 20165 14059 20223 14065
rect 20165 14056 20177 14059
rect 20128 14028 20177 14056
rect 20128 14016 20134 14028
rect 20165 14025 20177 14028
rect 20211 14025 20223 14059
rect 20165 14019 20223 14025
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20901 14059 20959 14065
rect 20901 14025 20913 14059
rect 20947 14056 20959 14059
rect 20990 14056 20996 14068
rect 20947 14028 20996 14056
rect 20947 14025 20959 14028
rect 20901 14019 20959 14025
rect 20990 14016 20996 14028
rect 21048 14016 21054 14068
rect 22922 14016 22928 14068
rect 22980 14056 22986 14068
rect 22980 14028 26280 14056
rect 22980 14016 22986 14028
rect 14660 13960 20484 13988
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 14148 13892 14381 13920
rect 14148 13880 14154 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13889 14519 13923
rect 14568 13920 14596 13948
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 14568 13892 14657 13920
rect 14461 13883 14519 13889
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 16022 13880 16028 13932
rect 16080 13920 16086 13932
rect 16117 13923 16175 13929
rect 16117 13920 16129 13923
rect 16080 13892 16129 13920
rect 16080 13880 16086 13892
rect 16117 13889 16129 13892
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16853 13923 16911 13929
rect 16853 13889 16865 13923
rect 16899 13920 16911 13923
rect 17034 13920 17040 13932
rect 16899 13892 17040 13920
rect 16899 13889 16911 13892
rect 16853 13883 16911 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 18138 13920 18144 13932
rect 17359 13892 18144 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 18230 13880 18236 13932
rect 18288 13880 18294 13932
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13920 18475 13923
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18463 13892 18521 13920
rect 18463 13889 18475 13892
rect 18417 13883 18475 13889
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 13136 13824 13216 13852
rect 13136 13812 13142 13824
rect 13538 13812 13544 13864
rect 13596 13812 13602 13864
rect 13648 13852 13676 13880
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13648 13824 13921 13852
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 14016 13852 14044 13880
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14016 13824 14565 13852
rect 13909 13815 13967 13821
rect 14553 13821 14565 13824
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 17402 13812 17408 13864
rect 17460 13812 17466 13864
rect 18524 13852 18552 13883
rect 18690 13880 18696 13932
rect 18748 13880 18754 13932
rect 19334 13852 19340 13864
rect 18524 13824 19340 13852
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13821 20407 13855
rect 20456 13852 20484 13960
rect 20622 13948 20628 14000
rect 20680 13988 20686 14000
rect 20680 13960 22600 13988
rect 20680 13948 20686 13960
rect 20990 13880 20996 13932
rect 21048 13880 21054 13932
rect 22572 13929 22600 13960
rect 23474 13948 23480 14000
rect 23532 13948 23538 14000
rect 26252 13988 26280 14028
rect 28902 14016 28908 14068
rect 28960 14016 28966 14068
rect 29089 13991 29147 13997
rect 29089 13988 29101 13991
rect 26252 13960 29101 13988
rect 29089 13957 29101 13960
rect 29135 13957 29147 13991
rect 29089 13951 29147 13957
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 20456 13824 21956 13852
rect 20349 13815 20407 13821
rect 13817 13787 13875 13793
rect 13817 13784 13829 13787
rect 13004 13756 13829 13784
rect 11020 13744 11026 13756
rect 13817 13753 13829 13756
rect 13863 13753 13875 13787
rect 13817 13747 13875 13753
rect 14642 13744 14648 13796
rect 14700 13784 14706 13796
rect 19426 13784 19432 13796
rect 14700 13756 19432 13784
rect 14700 13744 14706 13756
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 19794 13744 19800 13796
rect 19852 13784 19858 13796
rect 19978 13784 19984 13796
rect 19852 13756 19984 13784
rect 19852 13744 19858 13756
rect 19978 13744 19984 13756
rect 20036 13784 20042 13796
rect 20364 13784 20392 13815
rect 21928 13784 21956 13824
rect 22002 13812 22008 13864
rect 22060 13812 22066 13864
rect 22112 13852 22140 13883
rect 26050 13880 26056 13932
rect 26108 13880 26114 13932
rect 28810 13880 28816 13932
rect 28868 13920 28874 13932
rect 28997 13923 29055 13929
rect 28997 13920 29009 13923
rect 28868 13892 29009 13920
rect 28868 13880 28874 13892
rect 28997 13889 29009 13892
rect 29043 13889 29055 13923
rect 28997 13883 29055 13889
rect 29270 13880 29276 13932
rect 29328 13880 29334 13932
rect 23198 13852 23204 13864
rect 22112 13824 23204 13852
rect 23198 13812 23204 13824
rect 23256 13852 23262 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23256 13824 24593 13852
rect 23256 13812 23262 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 24673 13855 24731 13861
rect 24673 13821 24685 13855
rect 24719 13821 24731 13855
rect 24673 13815 24731 13821
rect 22278 13784 22284 13796
rect 20036 13756 20484 13784
rect 21928 13756 22284 13784
rect 20036 13744 20042 13756
rect 7156 13688 8064 13716
rect 7156 13676 7162 13688
rect 9030 13676 9036 13728
rect 9088 13676 9094 13728
rect 9769 13719 9827 13725
rect 9769 13685 9781 13719
rect 9815 13716 9827 13719
rect 10502 13716 10508 13728
rect 9815 13688 10508 13716
rect 9815 13685 9827 13688
rect 9769 13679 9827 13685
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 11238 13676 11244 13728
rect 11296 13676 11302 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12618 13716 12624 13728
rect 11664 13688 12624 13716
rect 11664 13676 11670 13688
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12802 13676 12808 13728
rect 12860 13676 12866 13728
rect 15654 13676 15660 13728
rect 15712 13676 15718 13728
rect 16758 13676 16764 13728
rect 16816 13676 16822 13728
rect 20456 13716 20484 13756
rect 22278 13744 22284 13756
rect 22336 13744 22342 13796
rect 22094 13716 22100 13728
rect 20456 13688 22100 13716
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 22373 13719 22431 13725
rect 22373 13685 22385 13719
rect 22419 13716 22431 13719
rect 22814 13719 22872 13725
rect 22814 13716 22826 13719
rect 22419 13688 22826 13716
rect 22419 13685 22431 13688
rect 22373 13679 22431 13685
rect 22814 13685 22826 13688
rect 22860 13685 22872 13719
rect 24688 13716 24716 13815
rect 24946 13812 24952 13864
rect 25004 13812 25010 13864
rect 27154 13812 27160 13864
rect 27212 13812 27218 13864
rect 27522 13744 27528 13796
rect 27580 13744 27586 13796
rect 25130 13716 25136 13728
rect 24688 13688 25136 13716
rect 22814 13679 22872 13685
rect 25130 13676 25136 13688
rect 25188 13676 25194 13728
rect 26418 13676 26424 13728
rect 26476 13676 26482 13728
rect 27617 13719 27675 13725
rect 27617 13685 27629 13719
rect 27663 13716 27675 13719
rect 27890 13716 27896 13728
rect 27663 13688 27896 13716
rect 27663 13685 27675 13688
rect 27617 13679 27675 13685
rect 27890 13676 27896 13688
rect 27948 13676 27954 13728
rect 1104 13626 29716 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 29716 13626
rect 1104 13552 29716 13574
rect 3786 13472 3792 13524
rect 3844 13472 3850 13524
rect 11330 13472 11336 13524
rect 11388 13512 11394 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11388 13484 11621 13512
rect 11388 13472 11394 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 11624 13444 11652 13475
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11848 13484 12081 13512
rect 11848 13472 11854 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 20438 13512 20444 13524
rect 19484 13484 20444 13512
rect 19484 13472 19490 13484
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 23474 13472 23480 13524
rect 23532 13472 23538 13524
rect 26050 13472 26056 13524
rect 26108 13512 26114 13524
rect 26329 13515 26387 13521
rect 26329 13512 26341 13515
rect 26108 13484 26341 13512
rect 26108 13472 26114 13484
rect 26329 13481 26341 13484
rect 26375 13481 26387 13515
rect 26329 13475 26387 13481
rect 27154 13472 27160 13524
rect 27212 13512 27218 13524
rect 27525 13515 27583 13521
rect 27525 13512 27537 13515
rect 27212 13484 27537 13512
rect 27212 13472 27218 13484
rect 27525 13481 27537 13484
rect 27571 13481 27583 13515
rect 27525 13475 27583 13481
rect 11624 13416 12296 13444
rect 2590 13336 2596 13388
rect 2648 13336 2654 13388
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 4706 13376 4712 13388
rect 4479 13348 4712 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 11238 13376 11244 13388
rect 10520 13348 11244 13376
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 2498 13308 2504 13320
rect 2087 13280 2504 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13308 2743 13311
rect 3510 13308 3516 13320
rect 2731 13280 3516 13308
rect 2731 13277 2743 13280
rect 2685 13271 2743 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4249 13311 4307 13317
rect 4249 13308 4261 13311
rect 4120 13280 4261 13308
rect 4120 13268 4126 13280
rect 4249 13277 4261 13280
rect 4295 13308 4307 13311
rect 7190 13308 7196 13320
rect 4295 13280 7196 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7650 13268 7656 13320
rect 7708 13268 7714 13320
rect 7926 13268 7932 13320
rect 7984 13268 7990 13320
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 10520 13317 10548 13348
rect 11238 13336 11244 13348
rect 11296 13336 11302 13388
rect 11808 13348 12204 13376
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 8168 13280 8217 13308
rect 8168 13268 8174 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 10594 13268 10600 13320
rect 10652 13268 10658 13320
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 3068 13212 4169 13240
rect 2130 13132 2136 13184
rect 2188 13132 2194 13184
rect 3068 13181 3096 13212
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 4157 13203 4215 13209
rect 6270 13200 6276 13252
rect 6328 13200 6334 13252
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13240 6515 13243
rect 6546 13240 6552 13252
rect 6503 13212 6552 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 6546 13200 6552 13212
rect 6604 13200 6610 13252
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7340 13212 8156 13240
rect 7340 13200 7346 13212
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13141 3111 13175
rect 3053 13135 3111 13141
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13172 7527 13175
rect 7558 13172 7564 13184
rect 7515 13144 7564 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7558 13132 7564 13144
rect 7616 13132 7622 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 8128 13181 8156 13212
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 10796 13240 10824 13271
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11808 13317 11836 13348
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13308 11115 13311
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11103 13280 11805 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 12066 13308 12072 13320
rect 11931 13280 12072 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 12176 13317 12204 13348
rect 12268 13317 12296 13416
rect 12434 13404 12440 13456
rect 12492 13444 12498 13456
rect 12529 13447 12587 13453
rect 12529 13444 12541 13447
rect 12492 13416 12541 13444
rect 12492 13404 12498 13416
rect 12529 13413 12541 13416
rect 12575 13413 12587 13447
rect 12529 13407 12587 13413
rect 22002 13404 22008 13456
rect 22060 13444 22066 13456
rect 27614 13444 27620 13456
rect 22060 13416 23428 13444
rect 22060 13404 22066 13416
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 15013 13379 15071 13385
rect 15013 13376 15025 13379
rect 14332 13348 15025 13376
rect 14332 13336 14338 13348
rect 15013 13345 15025 13348
rect 15059 13345 15071 13379
rect 15013 13339 15071 13345
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15654 13376 15660 13388
rect 15335 13348 15660 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16022 13336 16028 13388
rect 16080 13376 16086 13388
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 16080 13348 17049 13376
rect 16080 13336 16086 13348
rect 17037 13345 17049 13348
rect 17083 13376 17095 13379
rect 18230 13376 18236 13388
rect 17083 13348 18236 13376
rect 17083 13345 17095 13348
rect 17037 13339 17095 13345
rect 18230 13336 18236 13348
rect 18288 13376 18294 13388
rect 18690 13376 18696 13388
rect 18288 13348 18696 13376
rect 18288 13336 18294 13348
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 12254 13311 12312 13317
rect 12254 13277 12266 13311
rect 12300 13277 12312 13311
rect 12254 13271 12312 13277
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 12860 13280 13277 13308
rect 12860 13268 12866 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13446 13268 13452 13320
rect 13504 13268 13510 13320
rect 17126 13268 17132 13320
rect 17184 13308 17190 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17184 13280 17693 13308
rect 17184 13268 17190 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 8536 13212 10824 13240
rect 8536 13200 8542 13212
rect 11606 13200 11612 13252
rect 11664 13200 11670 13252
rect 16758 13240 16764 13252
rect 16514 13212 16764 13240
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 17696 13240 17724 13271
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 20349 13311 20407 13317
rect 20349 13308 20361 13311
rect 19392 13280 20361 13308
rect 19392 13268 19398 13280
rect 20349 13277 20361 13280
rect 20395 13308 20407 13311
rect 20395 13280 20576 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20438 13240 20444 13252
rect 17696 13212 20444 13240
rect 20438 13200 20444 13212
rect 20496 13200 20502 13252
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7800 13144 7849 13172
rect 7800 13132 7806 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 7837 13135 7895 13141
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 9490 13172 9496 13184
rect 8159 13144 9496 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 9490 13132 9496 13144
rect 9548 13132 9554 13184
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 12952 13144 13645 13172
rect 12952 13132 12958 13144
rect 13633 13141 13645 13144
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 17678 13132 17684 13184
rect 17736 13172 17742 13184
rect 17773 13175 17831 13181
rect 17773 13172 17785 13175
rect 17736 13144 17785 13172
rect 17736 13132 17742 13144
rect 17773 13141 17785 13144
rect 17819 13141 17831 13175
rect 20548 13172 20576 13280
rect 20622 13268 20628 13320
rect 20680 13268 20686 13320
rect 23400 13317 23428 13416
rect 26160 13416 27620 13444
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 26160 13385 26188 13416
rect 27614 13404 27620 13416
rect 27672 13404 27678 13456
rect 26145 13379 26203 13385
rect 26145 13376 26157 13379
rect 25188 13348 26157 13376
rect 25188 13336 25194 13348
rect 26145 13345 26157 13348
rect 26191 13345 26203 13379
rect 26145 13339 26203 13345
rect 27890 13336 27896 13388
rect 27948 13336 27954 13388
rect 23385 13311 23443 13317
rect 23385 13277 23397 13311
rect 23431 13277 23443 13311
rect 23385 13271 23443 13277
rect 24121 13311 24179 13317
rect 24121 13277 24133 13311
rect 24167 13308 24179 13311
rect 25148 13308 25176 13336
rect 24167 13280 25176 13308
rect 24167 13277 24179 13280
rect 24121 13271 24179 13277
rect 26326 13268 26332 13320
rect 26384 13308 26390 13320
rect 26421 13311 26479 13317
rect 26421 13308 26433 13311
rect 26384 13280 26433 13308
rect 26384 13268 26390 13280
rect 26421 13277 26433 13280
rect 26467 13308 26479 13311
rect 26878 13308 26884 13320
rect 26467 13280 26884 13308
rect 26467 13277 26479 13280
rect 26421 13271 26479 13277
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 26973 13311 27031 13317
rect 26973 13277 26985 13311
rect 27019 13308 27031 13311
rect 27154 13308 27160 13320
rect 27019 13280 27160 13308
rect 27019 13277 27031 13280
rect 26973 13271 27031 13277
rect 27154 13268 27160 13280
rect 27212 13268 27218 13320
rect 27249 13311 27307 13317
rect 27249 13277 27261 13311
rect 27295 13308 27307 13311
rect 27295 13280 27568 13308
rect 27295 13277 27307 13280
rect 27249 13271 27307 13277
rect 20898 13200 20904 13252
rect 20956 13200 20962 13252
rect 21910 13200 21916 13252
rect 21968 13200 21974 13252
rect 24210 13200 24216 13252
rect 24268 13240 24274 13252
rect 24397 13243 24455 13249
rect 24397 13240 24409 13243
rect 24268 13212 24409 13240
rect 24268 13200 24274 13212
rect 24397 13209 24409 13212
rect 24443 13209 24455 13243
rect 24397 13203 24455 13209
rect 27062 13200 27068 13252
rect 27120 13240 27126 13252
rect 27540 13240 27568 13280
rect 27614 13268 27620 13320
rect 27672 13268 27678 13320
rect 27120 13212 27936 13240
rect 27120 13200 27126 13212
rect 20714 13172 20720 13184
rect 20548 13144 20720 13172
rect 17773 13135 17831 13141
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22370 13132 22376 13184
rect 22428 13132 22434 13184
rect 26602 13132 26608 13184
rect 26660 13172 26666 13184
rect 27157 13175 27215 13181
rect 27157 13172 27169 13175
rect 26660 13144 27169 13172
rect 26660 13132 26666 13144
rect 27157 13141 27169 13144
rect 27203 13172 27215 13175
rect 27246 13172 27252 13184
rect 27203 13144 27252 13172
rect 27203 13141 27215 13144
rect 27157 13135 27215 13141
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 27341 13175 27399 13181
rect 27341 13141 27353 13175
rect 27387 13172 27399 13175
rect 27706 13172 27712 13184
rect 27387 13144 27712 13172
rect 27387 13141 27399 13144
rect 27341 13135 27399 13141
rect 27706 13132 27712 13144
rect 27764 13132 27770 13184
rect 27908 13172 27936 13212
rect 28902 13200 28908 13252
rect 28960 13200 28966 13252
rect 29365 13175 29423 13181
rect 29365 13172 29377 13175
rect 27908 13144 29377 13172
rect 29365 13141 29377 13144
rect 29411 13141 29423 13175
rect 29365 13135 29423 13141
rect 1104 13082 29716 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 29716 13082
rect 1104 13008 29716 13030
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 3786 12968 3792 12980
rect 3568 12940 3792 12968
rect 3568 12928 3574 12940
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 5997 12971 6055 12977
rect 5997 12937 6009 12971
rect 6043 12937 6055 12971
rect 5997 12931 6055 12937
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 6822 12968 6828 12980
rect 6779 12940 6828 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 1946 12900 1952 12912
rect 1412 12872 1952 12900
rect 1412 12841 1440 12872
rect 1946 12860 1952 12872
rect 2004 12860 2010 12912
rect 2130 12860 2136 12912
rect 2188 12860 2194 12912
rect 4798 12900 4804 12912
rect 4264 12872 4804 12900
rect 1397 12835 1455 12841
rect 1397 12801 1409 12835
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4062 12832 4068 12844
rect 3927 12804 4068 12832
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4264 12841 4292 12872
rect 4798 12860 4804 12872
rect 4856 12860 4862 12912
rect 5534 12860 5540 12912
rect 5592 12860 5598 12912
rect 6012 12900 6040 12931
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7834 12968 7840 12980
rect 7760 12940 7840 12968
rect 6270 12900 6276 12912
rect 6012 12872 6276 12900
rect 6270 12860 6276 12872
rect 6328 12900 6334 12912
rect 6641 12903 6699 12909
rect 6641 12900 6653 12903
rect 6328 12872 6653 12900
rect 6328 12860 6334 12872
rect 6641 12869 6653 12872
rect 6687 12900 6699 12903
rect 6687 12872 7696 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 6546 12792 6552 12844
rect 6604 12792 6610 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 7190 12832 7196 12844
rect 6788 12804 7196 12832
rect 6788 12792 6794 12804
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7340 12804 7389 12832
rect 7340 12792 7346 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7377 12795 7435 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 3418 12724 3424 12776
rect 3476 12724 3482 12776
rect 3970 12724 3976 12776
rect 4028 12724 4034 12776
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5994 12764 6000 12776
rect 4571 12736 6000 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 7006 12764 7012 12776
rect 6963 12736 7012 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 4614 12588 4620 12640
rect 4672 12628 4678 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 4672 12600 6377 12628
rect 4672 12588 4678 12600
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 6365 12591 6423 12597
rect 7377 12631 7435 12637
rect 7377 12597 7389 12631
rect 7423 12628 7435 12631
rect 7484 12628 7512 12795
rect 7558 12792 7564 12844
rect 7616 12792 7622 12844
rect 7668 12696 7696 12872
rect 7760 12841 7788 12940
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7984 12940 8309 12968
rect 7984 12928 7990 12940
rect 8297 12937 8309 12940
rect 8343 12968 8355 12971
rect 9033 12971 9091 12977
rect 8343 12940 8616 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 8588 12900 8616 12940
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9079 12940 9873 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 10318 12968 10324 12980
rect 9861 12931 9919 12937
rect 9968 12940 10324 12968
rect 9309 12903 9367 12909
rect 9309 12900 9321 12903
rect 8588 12872 9321 12900
rect 7745 12835 7803 12841
rect 7745 12801 7757 12835
rect 7791 12801 7803 12835
rect 7745 12795 7803 12801
rect 7837 12835 7895 12841
rect 7837 12801 7849 12835
rect 7883 12832 7895 12835
rect 7926 12832 7932 12844
rect 7883 12804 7932 12832
rect 7883 12801 7895 12804
rect 7837 12795 7895 12801
rect 7760 12764 7788 12795
rect 7926 12792 7932 12804
rect 7984 12832 7990 12844
rect 8202 12832 8208 12844
rect 7984 12804 8208 12832
rect 7984 12792 7990 12804
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 7760 12736 8248 12764
rect 8220 12708 8248 12736
rect 7668 12668 8156 12696
rect 7650 12628 7656 12640
rect 7423 12600 7656 12628
rect 7423 12597 7435 12600
rect 7377 12591 7435 12597
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 7834 12588 7840 12640
rect 7892 12628 7898 12640
rect 8021 12631 8079 12637
rect 8021 12628 8033 12631
rect 7892 12600 8033 12628
rect 7892 12588 7898 12600
rect 8021 12597 8033 12600
rect 8067 12597 8079 12631
rect 8128 12628 8156 12668
rect 8202 12656 8208 12708
rect 8260 12656 8266 12708
rect 8496 12696 8524 12792
rect 8588 12773 8616 12872
rect 9309 12869 9321 12872
rect 9355 12869 9367 12903
rect 9309 12863 9367 12869
rect 9401 12903 9459 12909
rect 9401 12869 9413 12903
rect 9447 12900 9459 12903
rect 9968 12900 9996 12940
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 14568 12940 16160 12968
rect 9447 12872 9996 12900
rect 10045 12903 10103 12909
rect 9447 12869 9459 12872
rect 9401 12863 9459 12869
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10226 12900 10232 12912
rect 10091 12872 10232 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12801 8815 12835
rect 8757 12795 8815 12801
rect 8573 12767 8631 12773
rect 8573 12733 8585 12767
rect 8619 12733 8631 12767
rect 8772 12764 8800 12795
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9030 12832 9036 12844
rect 8904 12804 9036 12832
rect 8904 12792 8910 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 8938 12764 8944 12776
rect 8772 12736 8944 12764
rect 8573 12727 8631 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 9140 12696 9168 12795
rect 9490 12792 9496 12844
rect 9548 12792 9554 12844
rect 9766 12792 9772 12844
rect 9824 12792 9830 12844
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 9508 12764 9536 12792
rect 10152 12764 10180 12795
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11422 12832 11428 12844
rect 11287 12804 11428 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 14274 12792 14280 12844
rect 14332 12832 14338 12844
rect 14568 12841 14596 12940
rect 14826 12860 14832 12912
rect 14884 12860 14890 12912
rect 15838 12860 15844 12912
rect 15896 12860 15902 12912
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 14332 12804 14565 12832
rect 14332 12792 14338 12804
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 16132 12832 16160 12940
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 17920 12940 18429 12968
rect 17920 12928 17926 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 19702 12968 19708 12980
rect 18417 12931 18475 12937
rect 18616 12940 19708 12968
rect 17678 12860 17684 12912
rect 17736 12860 17742 12912
rect 18616 12841 18644 12940
rect 19702 12928 19708 12940
rect 19760 12968 19766 12980
rect 20622 12968 20628 12980
rect 19760 12940 20628 12968
rect 19760 12928 19766 12940
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 20898 12928 20904 12980
rect 20956 12928 20962 12980
rect 21910 12928 21916 12980
rect 21968 12928 21974 12980
rect 24946 12928 24952 12980
rect 25004 12968 25010 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 25004 12940 25053 12968
rect 25004 12928 25010 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 26418 12968 26424 12980
rect 25041 12931 25099 12937
rect 25424 12940 26424 12968
rect 20533 12903 20591 12909
rect 20533 12900 20545 12903
rect 20102 12872 20545 12900
rect 20533 12869 20545 12872
rect 20579 12869 20591 12903
rect 20533 12863 20591 12869
rect 21266 12860 21272 12912
rect 21324 12860 21330 12912
rect 21361 12903 21419 12909
rect 21361 12869 21373 12903
rect 21407 12900 21419 12903
rect 22370 12900 22376 12912
rect 21407 12872 22376 12900
rect 21407 12869 21419 12872
rect 21361 12863 21419 12869
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16132 12804 16681 12832
rect 14553 12795 14611 12801
rect 16669 12801 16681 12804
rect 16715 12801 16727 12835
rect 16669 12795 16727 12801
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 20496 12804 20637 12832
rect 20496 12792 20502 12804
rect 20625 12801 20637 12804
rect 20671 12832 20683 12835
rect 20990 12832 20996 12844
rect 20671 12804 20996 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 20990 12792 20996 12804
rect 21048 12832 21054 12844
rect 22002 12832 22008 12844
rect 21048 12804 22008 12832
rect 21048 12792 21054 12804
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 25424 12841 25452 12940
rect 26418 12928 26424 12940
rect 26476 12968 26482 12980
rect 27154 12968 27160 12980
rect 26476 12940 27160 12968
rect 26476 12928 26482 12940
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 27522 12928 27528 12980
rect 27580 12928 27586 12980
rect 28813 12971 28871 12977
rect 28813 12937 28825 12971
rect 28859 12968 28871 12971
rect 28902 12968 28908 12980
rect 28859 12940 28908 12968
rect 28859 12937 28871 12940
rect 28813 12931 28871 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 27617 12903 27675 12909
rect 27617 12900 27629 12903
rect 25884 12872 27629 12900
rect 25884 12841 25912 12872
rect 27617 12869 27629 12872
rect 27663 12869 27675 12903
rect 27617 12863 27675 12869
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 26602 12792 26608 12844
rect 26660 12792 26666 12844
rect 26789 12835 26847 12841
rect 26789 12801 26801 12835
rect 26835 12801 26847 12835
rect 26789 12795 26847 12801
rect 9508 12736 10180 12764
rect 10410 12724 10416 12776
rect 10468 12764 10474 12776
rect 10468 12736 16436 12764
rect 10468 12724 10474 12736
rect 8496 12668 9168 12696
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 10226 12696 10232 12708
rect 9723 12668 10232 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 10226 12656 10232 12668
rect 10284 12656 10290 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 11514 12696 11520 12708
rect 10836 12668 11520 12696
rect 10836 12656 10842 12668
rect 11514 12656 11520 12668
rect 11572 12696 11578 12708
rect 13078 12696 13084 12708
rect 11572 12668 13084 12696
rect 11572 12656 11578 12668
rect 13078 12656 13084 12668
rect 13136 12696 13142 12708
rect 13630 12696 13636 12708
rect 13136 12668 13636 12696
rect 13136 12656 13142 12668
rect 13630 12656 13636 12668
rect 13688 12656 13694 12708
rect 8938 12628 8944 12640
rect 8128 12600 8944 12628
rect 8021 12591 8079 12597
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 10042 12588 10048 12640
rect 10100 12588 10106 12640
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 11146 12588 11152 12640
rect 11204 12588 11210 12640
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 16301 12631 16359 12637
rect 16301 12628 16313 12631
rect 14976 12600 16313 12628
rect 14976 12588 14982 12600
rect 16301 12597 16313 12600
rect 16347 12597 16359 12631
rect 16408 12628 16436 12736
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 18874 12724 18880 12776
rect 18932 12724 18938 12776
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 22094 12764 22100 12776
rect 21591 12736 22100 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 22094 12724 22100 12736
rect 22152 12764 22158 12776
rect 23658 12764 23664 12776
rect 22152 12736 23664 12764
rect 22152 12724 22158 12736
rect 23658 12724 23664 12736
rect 23716 12724 23722 12776
rect 25501 12767 25559 12773
rect 25501 12733 25513 12767
rect 25547 12764 25559 12767
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25547 12736 26065 12764
rect 25547 12733 25559 12736
rect 25501 12727 25559 12733
rect 26053 12733 26065 12736
rect 26099 12764 26111 12767
rect 26697 12767 26755 12773
rect 26697 12764 26709 12767
rect 26099 12736 26709 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 26697 12733 26709 12736
rect 26743 12733 26755 12767
rect 26804 12764 26832 12795
rect 27062 12792 27068 12844
rect 27120 12792 27126 12844
rect 27154 12792 27160 12844
rect 27212 12792 27218 12844
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 27430 12832 27436 12844
rect 27304 12804 27436 12832
rect 27304 12792 27310 12804
rect 27430 12792 27436 12804
rect 27488 12832 27494 12844
rect 27801 12835 27859 12841
rect 27801 12832 27813 12835
rect 27488 12804 27813 12832
rect 27488 12792 27494 12804
rect 27801 12801 27813 12804
rect 27847 12801 27859 12835
rect 27801 12795 27859 12801
rect 27982 12792 27988 12844
rect 28040 12792 28046 12844
rect 28810 12792 28816 12844
rect 28868 12832 28874 12844
rect 28905 12835 28963 12841
rect 28905 12832 28917 12835
rect 28868 12804 28917 12832
rect 28868 12792 28874 12804
rect 28905 12801 28917 12804
rect 28951 12801 28963 12835
rect 28905 12795 28963 12801
rect 29270 12792 29276 12844
rect 29328 12792 29334 12844
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 26804 12736 27353 12764
rect 26697 12727 26755 12733
rect 27341 12733 27353 12736
rect 27387 12764 27399 12767
rect 27706 12764 27712 12776
rect 27387 12736 27712 12764
rect 27387 12733 27399 12736
rect 27341 12727 27399 12733
rect 27706 12724 27712 12736
rect 27764 12764 27770 12776
rect 28000 12764 28028 12792
rect 27764 12736 28028 12764
rect 27764 12724 27770 12736
rect 29089 12699 29147 12705
rect 29089 12696 29101 12699
rect 19904 12668 29101 12696
rect 19904 12628 19932 12668
rect 29089 12665 29101 12668
rect 29135 12665 29147 12699
rect 29089 12659 29147 12665
rect 16408 12600 19932 12628
rect 16301 12591 16359 12597
rect 20346 12588 20352 12640
rect 20404 12588 20410 12640
rect 25682 12588 25688 12640
rect 25740 12588 25746 12640
rect 1104 12538 29716 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 29716 12538
rect 1104 12464 29716 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1728 12396 1869 12424
rect 1728 12384 1734 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 2498 12384 2504 12436
rect 2556 12424 2562 12436
rect 5261 12427 5319 12433
rect 2556 12396 5212 12424
rect 2556 12384 2562 12396
rect 3326 12356 3332 12368
rect 2516 12328 3332 12356
rect 2516 12297 2544 12328
rect 3326 12316 3332 12328
rect 3384 12356 3390 12368
rect 4706 12356 4712 12368
rect 3384 12328 4712 12356
rect 3384 12316 3390 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 5184 12356 5212 12396
rect 5261 12393 5273 12427
rect 5307 12424 5319 12427
rect 5534 12424 5540 12436
rect 5307 12396 5540 12424
rect 5307 12393 5319 12396
rect 5261 12387 5319 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 5994 12384 6000 12436
rect 6052 12384 6058 12436
rect 6181 12427 6239 12433
rect 6181 12393 6193 12427
rect 6227 12424 6239 12427
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6227 12396 6561 12424
rect 6227 12393 6239 12396
rect 6181 12387 6239 12393
rect 6549 12393 6561 12396
rect 6595 12424 6607 12427
rect 6638 12424 6644 12436
rect 6595 12396 6644 12424
rect 6595 12393 6607 12396
rect 6549 12387 6607 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 7466 12424 7472 12436
rect 7340 12396 7472 12424
rect 7340 12384 7346 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 7650 12384 7656 12436
rect 7708 12384 7714 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 8812 12396 9597 12424
rect 8812 12384 8818 12396
rect 9585 12393 9597 12396
rect 9631 12393 9643 12427
rect 9585 12387 9643 12393
rect 10042 12384 10048 12436
rect 10100 12384 10106 12436
rect 10152 12396 10364 12424
rect 5442 12356 5448 12368
rect 5184 12328 5448 12356
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 3789 12291 3847 12297
rect 3789 12257 3801 12291
rect 3835 12288 3847 12291
rect 3970 12288 3976 12300
rect 3835 12260 3976 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 4062 12248 4068 12300
rect 4120 12248 4126 12300
rect 842 12180 848 12232
rect 900 12220 906 12232
rect 1489 12223 1547 12229
rect 1489 12220 1501 12223
rect 900 12192 1501 12220
rect 900 12180 906 12192
rect 1489 12189 1501 12192
rect 1535 12189 1547 12223
rect 1489 12183 1547 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3142 12220 3148 12232
rect 2363 12192 3148 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3142 12180 3148 12192
rect 3200 12220 3206 12232
rect 3418 12220 3424 12232
rect 3200 12192 3424 12220
rect 3200 12180 3206 12192
rect 3418 12180 3424 12192
rect 3476 12220 3482 12232
rect 5184 12229 5212 12328
rect 5442 12316 5448 12328
rect 5500 12316 5506 12368
rect 10152 12356 10180 12396
rect 6656 12328 10180 12356
rect 10229 12359 10287 12365
rect 6546 12248 6552 12300
rect 6604 12288 6610 12300
rect 6656 12288 6684 12328
rect 10229 12325 10241 12359
rect 10275 12325 10287 12359
rect 10336 12356 10364 12396
rect 10502 12384 10508 12436
rect 10560 12384 10566 12436
rect 11054 12384 11060 12436
rect 11112 12424 11118 12436
rect 11238 12424 11244 12436
rect 11112 12396 11244 12424
rect 11112 12384 11118 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 14461 12427 14519 12433
rect 14461 12393 14473 12427
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 14645 12427 14703 12433
rect 14645 12393 14657 12427
rect 14691 12424 14703 12427
rect 14826 12424 14832 12436
rect 14691 12396 14832 12424
rect 14691 12393 14703 12396
rect 14645 12387 14703 12393
rect 13262 12356 13268 12368
rect 10336 12328 13268 12356
rect 10229 12319 10287 12325
rect 6604 12260 6684 12288
rect 6604 12248 6610 12260
rect 4157 12223 4215 12229
rect 4157 12220 4169 12223
rect 3476 12192 4169 12220
rect 3476 12180 3482 12192
rect 4157 12189 4169 12192
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 6086 12180 6092 12232
rect 6144 12220 6150 12232
rect 6144 12189 6208 12220
rect 6144 12180 6147 12189
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 1946 12152 1952 12164
rect 1719 12124 1952 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 1946 12112 1952 12124
rect 2004 12112 2010 12164
rect 6135 12155 6147 12180
rect 6181 12158 6208 12189
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 6656 12229 6684 12260
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 7926 12288 7932 12300
rect 7883 12260 7932 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 10244 12288 10272 12319
rect 13262 12316 13268 12328
rect 13320 12356 13326 12368
rect 14093 12359 14151 12365
rect 14093 12356 14105 12359
rect 13320 12328 14105 12356
rect 13320 12316 13326 12328
rect 14093 12325 14105 12328
rect 14139 12325 14151 12359
rect 14476 12356 14504 12387
rect 14826 12384 14832 12396
rect 14884 12384 14890 12436
rect 15749 12427 15807 12433
rect 15749 12393 15761 12427
rect 15795 12424 15807 12427
rect 15838 12424 15844 12436
rect 15795 12396 15844 12424
rect 15795 12393 15807 12396
rect 15749 12387 15807 12393
rect 15838 12384 15844 12396
rect 15896 12384 15902 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 17000 12396 17233 12424
rect 17000 12384 17006 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 17221 12387 17279 12393
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18932 12396 19257 12424
rect 18932 12384 18938 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 27157 12427 27215 12433
rect 27157 12393 27169 12427
rect 27203 12424 27215 12427
rect 27430 12424 27436 12436
rect 27203 12396 27436 12424
rect 27203 12393 27215 12396
rect 27157 12387 27215 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 15105 12359 15163 12365
rect 15105 12356 15117 12359
rect 14476 12328 15117 12356
rect 14093 12319 14151 12325
rect 15105 12325 15117 12328
rect 15151 12325 15163 12359
rect 15105 12319 15163 12325
rect 9640 12260 9812 12288
rect 9640 12248 9646 12260
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 6328 12192 6469 12220
rect 6328 12180 6334 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7742 12220 7748 12232
rect 7616 12192 7748 12220
rect 7616 12180 7622 12192
rect 7742 12180 7748 12192
rect 7800 12180 7806 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8205 12223 8263 12229
rect 8205 12220 8217 12223
rect 8168 12192 8217 12220
rect 8168 12180 8174 12192
rect 8205 12189 8217 12192
rect 8251 12189 8263 12223
rect 8205 12183 8263 12189
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8352 12192 8401 12220
rect 8352 12180 8358 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 9674 12220 9680 12232
rect 8389 12183 8447 12189
rect 8496 12192 9680 12220
rect 6181 12155 6193 12158
rect 6135 12149 6193 12155
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 8496 12152 8524 12192
rect 9674 12180 9680 12192
rect 9732 12180 9738 12232
rect 9784 12229 9812 12260
rect 9876 12260 10272 12288
rect 10612 12260 11468 12288
rect 9876 12229 9904 12260
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10413 12223 10471 12229
rect 10413 12220 10425 12223
rect 10284 12192 10425 12220
rect 10284 12180 10290 12192
rect 10413 12189 10425 12192
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 6420 12124 8524 12152
rect 6420 12112 6426 12124
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 10612 12152 10640 12260
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 10870 12220 10876 12232
rect 10827 12192 10876 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 8996 12124 10640 12152
rect 8996 12112 9002 12124
rect 10686 12112 10692 12164
rect 10744 12112 10750 12164
rect 2222 12044 2228 12096
rect 2280 12044 2286 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8113 12087 8171 12093
rect 8113 12084 8125 12087
rect 7892 12056 8125 12084
rect 7892 12044 7898 12056
rect 8113 12053 8125 12056
rect 8159 12053 8171 12087
rect 8113 12047 8171 12053
rect 8294 12044 8300 12096
rect 8352 12044 8358 12096
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 10796 12084 10824 12183
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11072 12229 11100 12260
rect 11057 12223 11115 12229
rect 11057 12189 11069 12223
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 11146 12180 11152 12232
rect 11204 12180 11210 12232
rect 11440 12229 11468 12260
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 15746 12288 15752 12300
rect 11756 12260 15752 12288
rect 11756 12248 11762 12260
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 16206 12248 16212 12300
rect 16264 12288 16270 12300
rect 16390 12288 16396 12300
rect 16264 12260 16396 12288
rect 16264 12248 16270 12260
rect 16390 12248 16396 12260
rect 16448 12288 16454 12300
rect 17773 12291 17831 12297
rect 17773 12288 17785 12291
rect 16448 12260 17785 12288
rect 16448 12248 16454 12260
rect 17773 12257 17785 12260
rect 17819 12288 17831 12291
rect 19889 12291 19947 12297
rect 19889 12288 19901 12291
rect 17819 12260 19901 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 19889 12257 19901 12260
rect 19935 12288 19947 12291
rect 19978 12288 19984 12300
rect 19935 12260 19984 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 19978 12248 19984 12260
rect 20036 12248 20042 12300
rect 22373 12291 22431 12297
rect 22373 12257 22385 12291
rect 22419 12288 22431 12291
rect 23109 12291 23167 12297
rect 23109 12288 23121 12291
rect 22419 12260 23121 12288
rect 22419 12257 22431 12260
rect 22373 12251 22431 12257
rect 23109 12257 23121 12260
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23658 12248 23664 12300
rect 23716 12288 23722 12300
rect 24949 12291 25007 12297
rect 24949 12288 24961 12291
rect 23716 12260 24961 12288
rect 23716 12248 23722 12260
rect 24949 12257 24961 12260
rect 24995 12257 25007 12291
rect 24949 12251 25007 12257
rect 25682 12248 25688 12300
rect 25740 12248 25746 12300
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 12894 12180 12900 12232
rect 12952 12180 12958 12232
rect 12986 12180 12992 12232
rect 13044 12180 13050 12232
rect 13078 12180 13084 12232
rect 13136 12180 13142 12232
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12220 13323 12223
rect 13538 12220 13544 12232
rect 13311 12192 13544 12220
rect 13311 12189 13323 12192
rect 13265 12183 13323 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 15841 12223 15899 12229
rect 15841 12189 15853 12223
rect 15887 12220 15899 12223
rect 16666 12220 16672 12232
rect 15887 12192 16672 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16666 12180 16672 12192
rect 16724 12220 16730 12232
rect 17034 12220 17040 12232
rect 16724 12192 17040 12220
rect 16724 12180 16730 12192
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 19702 12180 19708 12232
rect 19760 12220 19766 12232
rect 20346 12220 20352 12232
rect 19760 12192 20352 12220
rect 19760 12180 19766 12192
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 21634 12220 21640 12232
rect 20772 12192 21640 12220
rect 20772 12180 20778 12192
rect 21634 12180 21640 12192
rect 21692 12220 21698 12232
rect 21821 12223 21879 12229
rect 21821 12220 21833 12223
rect 21692 12192 21833 12220
rect 21692 12180 21698 12192
rect 21821 12189 21833 12192
rect 21867 12189 21879 12223
rect 21821 12183 21879 12189
rect 22002 12180 22008 12232
rect 22060 12180 22066 12232
rect 22278 12180 22284 12232
rect 22336 12180 22342 12232
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 22830 12180 22836 12232
rect 22888 12220 22894 12232
rect 23198 12220 23204 12232
rect 22888 12192 23204 12220
rect 22888 12180 22894 12192
rect 23198 12180 23204 12192
rect 23256 12180 23262 12232
rect 25130 12180 25136 12232
rect 25188 12220 25194 12232
rect 25409 12223 25467 12229
rect 25409 12220 25421 12223
rect 25188 12192 25421 12220
rect 25188 12180 25194 12192
rect 25409 12189 25421 12192
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 26970 12180 26976 12232
rect 27028 12220 27034 12232
rect 27433 12223 27491 12229
rect 27433 12220 27445 12223
rect 27028 12192 27445 12220
rect 27028 12180 27034 12192
rect 27433 12189 27445 12192
rect 27479 12220 27491 12223
rect 28902 12220 28908 12232
rect 27479 12192 28908 12220
rect 27479 12189 27491 12192
rect 27433 12183 27491 12189
rect 28902 12180 28908 12192
rect 28960 12180 28966 12232
rect 10965 12155 11023 12161
rect 10965 12121 10977 12155
rect 11011 12152 11023 12155
rect 11330 12152 11336 12164
rect 11011 12124 11336 12152
rect 11011 12121 11023 12124
rect 10965 12115 11023 12121
rect 11330 12112 11336 12124
rect 11388 12112 11394 12164
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14737 12155 14795 12161
rect 14737 12152 14749 12155
rect 14240 12124 14749 12152
rect 14240 12112 14246 12124
rect 14737 12121 14749 12124
rect 14783 12121 14795 12155
rect 14737 12115 14795 12121
rect 21913 12155 21971 12161
rect 21913 12121 21925 12155
rect 21959 12152 21971 12155
rect 22480 12152 22508 12180
rect 24765 12155 24823 12161
rect 24765 12152 24777 12155
rect 21959 12124 22508 12152
rect 23584 12124 24777 12152
rect 21959 12121 21971 12124
rect 21913 12115 21971 12121
rect 9088 12056 10824 12084
rect 9088 12044 9094 12056
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 13998 12084 14004 12096
rect 13872 12056 14004 12084
rect 13872 12044 13878 12056
rect 13998 12044 14004 12056
rect 14056 12084 14062 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14056 12056 14473 12084
rect 14056 12044 14062 12056
rect 14461 12053 14473 12056
rect 14507 12084 14519 12087
rect 14550 12084 14556 12096
rect 14507 12056 14556 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 17589 12087 17647 12093
rect 17589 12084 17601 12087
rect 17552 12056 17601 12084
rect 17552 12044 17558 12056
rect 17589 12053 17601 12056
rect 17635 12053 17647 12087
rect 17589 12047 17647 12053
rect 17681 12087 17739 12093
rect 17681 12053 17693 12087
rect 17727 12084 17739 12087
rect 17862 12084 17868 12096
rect 17727 12056 17868 12084
rect 17727 12053 17739 12056
rect 17681 12047 17739 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 19518 12044 19524 12096
rect 19576 12084 19582 12096
rect 23584 12093 23612 12124
rect 24765 12121 24777 12124
rect 24811 12121 24823 12155
rect 27341 12155 27399 12161
rect 27341 12152 27353 12155
rect 26910 12124 27353 12152
rect 24765 12115 24823 12121
rect 27341 12121 27353 12124
rect 27387 12121 27399 12155
rect 27341 12115 27399 12121
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19576 12056 19625 12084
rect 19576 12044 19582 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 19613 12047 19671 12053
rect 23569 12087 23627 12093
rect 23569 12053 23581 12087
rect 23615 12053 23627 12087
rect 23569 12047 23627 12053
rect 23934 12044 23940 12096
rect 23992 12084 23998 12096
rect 24397 12087 24455 12093
rect 24397 12084 24409 12087
rect 23992 12056 24409 12084
rect 23992 12044 23998 12056
rect 24397 12053 24409 12056
rect 24443 12053 24455 12087
rect 24397 12047 24455 12053
rect 24486 12044 24492 12096
rect 24544 12084 24550 12096
rect 24857 12087 24915 12093
rect 24857 12084 24869 12087
rect 24544 12056 24869 12084
rect 24544 12044 24550 12056
rect 24857 12053 24869 12056
rect 24903 12053 24915 12087
rect 24857 12047 24915 12053
rect 1104 11994 29716 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 29716 11994
rect 1104 11920 29716 11942
rect 5537 11883 5595 11889
rect 5537 11849 5549 11883
rect 5583 11880 5595 11883
rect 5626 11880 5632 11892
rect 5583 11852 5632 11880
rect 5583 11849 5595 11852
rect 5537 11843 5595 11849
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 7466 11880 7472 11892
rect 7392 11852 7472 11880
rect 4062 11772 4068 11824
rect 4120 11812 4126 11824
rect 4798 11812 4804 11824
rect 4120 11784 4804 11812
rect 4120 11772 4126 11784
rect 4798 11772 4804 11784
rect 4856 11812 4862 11824
rect 5261 11815 5319 11821
rect 5261 11812 5273 11815
rect 4856 11784 5273 11812
rect 4856 11772 4862 11784
rect 5261 11781 5273 11784
rect 5307 11781 5319 11815
rect 5261 11775 5319 11781
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 7392 11753 7420 11852
rect 7466 11840 7472 11852
rect 7524 11880 7530 11892
rect 8294 11880 8300 11892
rect 7524 11852 8300 11880
rect 7524 11840 7530 11852
rect 8294 11840 8300 11852
rect 8352 11840 8358 11892
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9766 11880 9772 11892
rect 9631 11852 9772 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9766 11840 9772 11852
rect 9824 11880 9830 11892
rect 10502 11880 10508 11892
rect 9824 11852 10508 11880
rect 9824 11840 9830 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 10744 11852 11529 11880
rect 10744 11840 10750 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 17494 11840 17500 11892
rect 17552 11840 17558 11892
rect 27982 11880 27988 11892
rect 27356 11852 27988 11880
rect 7834 11772 7840 11824
rect 7892 11821 7898 11824
rect 7892 11815 7920 11821
rect 7908 11781 7920 11815
rect 7892 11775 7920 11781
rect 7892 11772 7898 11775
rect 8846 11772 8852 11824
rect 8904 11812 8910 11824
rect 8904 11784 9444 11812
rect 8904 11772 8910 11784
rect 9416 11756 9444 11784
rect 10134 11772 10140 11824
rect 10192 11812 10198 11824
rect 12437 11815 12495 11821
rect 10192 11784 12204 11812
rect 10192 11772 10198 11784
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 7377 11747 7435 11753
rect 5399 11716 7236 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 5184 11676 5212 11707
rect 5184 11648 5396 11676
rect 5368 11620 5396 11648
rect 7208 11620 7236 11716
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7616 11716 8125 11744
rect 7616 11704 7622 11716
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 9180 11716 9229 11744
rect 9180 11704 9186 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 9398 11704 9404 11756
rect 9456 11704 9462 11756
rect 10502 11704 10508 11756
rect 10560 11704 10566 11756
rect 10594 11704 10600 11756
rect 10652 11744 10658 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10652 11716 10701 11744
rect 10652 11704 10658 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10781 11747 10839 11753
rect 10781 11713 10793 11747
rect 10827 11713 10839 11747
rect 10781 11707 10839 11713
rect 10873 11750 10931 11753
rect 10962 11750 10968 11756
rect 10873 11747 10968 11750
rect 10873 11713 10885 11747
rect 10919 11722 10968 11747
rect 10919 11713 10931 11722
rect 10873 11707 10931 11713
rect 7650 11636 7656 11688
rect 7708 11636 7714 11688
rect 7742 11636 7748 11688
rect 7800 11636 7806 11688
rect 9858 11676 9864 11688
rect 7852 11648 9864 11676
rect 5350 11568 5356 11620
rect 5408 11568 5414 11620
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 7852 11608 7880 11648
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 7248 11580 7880 11608
rect 7248 11568 7254 11580
rect 8018 11568 8024 11620
rect 8076 11568 8082 11620
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9306 11608 9312 11620
rect 8996 11580 9312 11608
rect 8996 11568 9002 11580
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 10686 11608 10692 11620
rect 9732 11580 10692 11608
rect 9732 11568 9738 11580
rect 10686 11568 10692 11580
rect 10744 11568 10750 11620
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 6270 11540 6276 11552
rect 3476 11512 6276 11540
rect 3476 11500 3482 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 10796 11540 10824 11707
rect 10962 11704 10968 11722
rect 11020 11704 11026 11756
rect 11698 11753 11704 11756
rect 11696 11744 11704 11753
rect 11659 11716 11704 11744
rect 11696 11707 11704 11716
rect 11698 11704 11704 11707
rect 11756 11704 11762 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 11974 11744 11980 11756
rect 11931 11716 11980 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 11057 11611 11115 11617
rect 11057 11577 11069 11611
rect 11103 11608 11115 11611
rect 11238 11608 11244 11620
rect 11103 11580 11244 11608
rect 11103 11577 11115 11580
rect 11057 11571 11115 11577
rect 11238 11568 11244 11580
rect 11296 11568 11302 11620
rect 11808 11608 11836 11707
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12176 11753 12204 11784
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 14001 11815 14059 11821
rect 12483 11784 13032 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 13004 11756 13032 11784
rect 14001 11781 14013 11815
rect 14047 11812 14059 11815
rect 14047 11784 14228 11812
rect 14047 11781 14059 11784
rect 14001 11775 14059 11781
rect 14200 11756 14228 11784
rect 14550 11772 14556 11824
rect 14608 11772 14614 11824
rect 16482 11772 16488 11824
rect 16540 11812 16546 11824
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 16540 11784 21833 11812
rect 16540 11772 16546 11784
rect 21821 11781 21833 11784
rect 21867 11812 21879 11815
rect 24210 11812 24216 11824
rect 21867 11784 24216 11812
rect 21867 11781 21879 11784
rect 21821 11775 21879 11781
rect 24210 11772 24216 11784
rect 24268 11772 24274 11824
rect 25685 11815 25743 11821
rect 25685 11812 25697 11815
rect 25162 11784 25697 11812
rect 25685 11781 25697 11784
rect 25731 11781 25743 11815
rect 25685 11775 25743 11781
rect 12068 11747 12126 11753
rect 12068 11713 12080 11747
rect 12114 11713 12126 11747
rect 12068 11707 12126 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12083 11676 12111 11707
rect 12894 11704 12900 11756
rect 12952 11704 12958 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13173 11747 13231 11753
rect 13173 11744 13185 11747
rect 13044 11716 13185 11744
rect 13044 11704 13050 11716
rect 13173 11713 13185 11716
rect 13219 11713 13231 11747
rect 13173 11707 13231 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13449 11747 13507 11753
rect 13449 11713 13461 11747
rect 13495 11713 13507 11747
rect 13449 11707 13507 11713
rect 12710 11676 12716 11688
rect 12083 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 12802 11636 12808 11688
rect 12860 11636 12866 11688
rect 13372 11676 13400 11707
rect 13004 11648 13400 11676
rect 13004 11608 13032 11648
rect 11808 11580 13032 11608
rect 12912 11552 12940 11580
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 8260 11512 10824 11540
rect 8260 11500 8266 11512
rect 12526 11500 12532 11552
rect 12584 11500 12590 11552
rect 12894 11500 12900 11552
rect 12952 11500 12958 11552
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13464 11540 13492 11707
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 13725 11747 13783 11753
rect 13725 11744 13737 11747
rect 13596 11716 13737 11744
rect 13596 11704 13602 11716
rect 13725 11713 13737 11716
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 13906 11704 13912 11756
rect 13964 11704 13970 11756
rect 14093 11747 14151 11753
rect 14093 11713 14105 11747
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 14108 11676 14136 11707
rect 14182 11704 14188 11756
rect 14240 11704 14246 11756
rect 14826 11704 14832 11756
rect 14884 11704 14890 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17310 11744 17316 11756
rect 17175 11716 17316 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 15028 11676 15056 11707
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 19058 11704 19064 11756
rect 19116 11704 19122 11756
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 20441 11747 20499 11753
rect 20441 11713 20453 11747
rect 20487 11744 20499 11747
rect 20487 11716 20668 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 20640 11688 20668 11716
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20772 11716 21005 11744
rect 20772 11704 20778 11716
rect 20993 11713 21005 11716
rect 21039 11744 21051 11747
rect 23385 11747 23443 11753
rect 23385 11744 23397 11747
rect 21039 11716 23397 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 23385 11713 23397 11716
rect 23431 11744 23443 11747
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23431 11716 23673 11744
rect 23431 11713 23443 11716
rect 23385 11707 23443 11713
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 25777 11747 25835 11753
rect 25777 11713 25789 11747
rect 25823 11744 25835 11747
rect 26418 11744 26424 11756
rect 25823 11716 26424 11744
rect 25823 11713 25835 11716
rect 25777 11707 25835 11713
rect 26418 11704 26424 11716
rect 26476 11744 26482 11756
rect 26878 11744 26884 11756
rect 26476 11716 26884 11744
rect 26476 11704 26482 11716
rect 26878 11704 26884 11716
rect 26936 11704 26942 11756
rect 27356 11753 27384 11852
rect 27982 11840 27988 11852
rect 28040 11840 28046 11892
rect 27433 11815 27491 11821
rect 27433 11781 27445 11815
rect 27479 11812 27491 11815
rect 27893 11815 27951 11821
rect 27893 11812 27905 11815
rect 27479 11784 27905 11812
rect 27479 11781 27491 11784
rect 27433 11775 27491 11781
rect 27893 11781 27905 11784
rect 27939 11781 27951 11815
rect 27893 11775 27951 11781
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11713 27399 11747
rect 27341 11707 27399 11713
rect 27522 11704 27528 11756
rect 27580 11704 27586 11756
rect 28994 11704 29000 11756
rect 29052 11704 29058 11756
rect 14108 11648 15056 11676
rect 13722 11568 13728 11620
rect 13780 11608 13786 11620
rect 14108 11608 14136 11648
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 20530 11636 20536 11688
rect 20588 11636 20594 11688
rect 20622 11636 20628 11688
rect 20680 11636 20686 11688
rect 20809 11679 20867 11685
rect 20809 11645 20821 11679
rect 20855 11676 20867 11679
rect 21266 11676 21272 11688
rect 20855 11648 21272 11676
rect 20855 11645 20867 11648
rect 20809 11639 20867 11645
rect 21266 11636 21272 11648
rect 21324 11636 21330 11688
rect 23934 11636 23940 11688
rect 23992 11636 23998 11688
rect 27614 11636 27620 11688
rect 27672 11636 27678 11688
rect 14921 11611 14979 11617
rect 14921 11608 14933 11611
rect 13780 11580 14136 11608
rect 14568 11580 14933 11608
rect 13780 11568 13786 11580
rect 14568 11549 14596 11580
rect 14921 11577 14933 11580
rect 14967 11577 14979 11611
rect 14921 11571 14979 11577
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 21910 11608 21916 11620
rect 15068 11580 21916 11608
rect 15068 11568 15074 11580
rect 21910 11568 21916 11580
rect 21968 11568 21974 11620
rect 23474 11608 23480 11620
rect 22066 11580 23480 11608
rect 13044 11512 13492 11540
rect 14553 11543 14611 11549
rect 13044 11500 13050 11512
rect 14553 11509 14565 11543
rect 14599 11509 14611 11543
rect 14553 11503 14611 11509
rect 14734 11500 14740 11552
rect 14792 11500 14798 11552
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19978 11540 19984 11552
rect 19291 11512 19984 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 21818 11500 21824 11552
rect 21876 11540 21882 11552
rect 22066 11540 22094 11580
rect 23474 11568 23480 11580
rect 23532 11568 23538 11620
rect 21876 11512 22094 11540
rect 21876 11500 21882 11512
rect 22370 11500 22376 11552
rect 22428 11540 22434 11552
rect 23014 11540 23020 11552
rect 22428 11512 23020 11540
rect 22428 11500 22434 11512
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 24486 11500 24492 11552
rect 24544 11540 24550 11552
rect 25409 11543 25467 11549
rect 25409 11540 25421 11543
rect 24544 11512 25421 11540
rect 24544 11500 24550 11512
rect 25409 11509 25421 11512
rect 25455 11509 25467 11543
rect 25409 11503 25467 11509
rect 28258 11500 28264 11552
rect 28316 11540 28322 11552
rect 29365 11543 29423 11549
rect 29365 11540 29377 11543
rect 28316 11512 29377 11540
rect 28316 11500 28322 11512
rect 29365 11509 29377 11512
rect 29411 11509 29423 11543
rect 29365 11503 29423 11509
rect 1104 11450 29716 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 29716 11450
rect 1104 11376 29716 11398
rect 1857 11339 1915 11345
rect 1857 11305 1869 11339
rect 1903 11336 1915 11339
rect 2222 11336 2228 11348
rect 1903 11308 2228 11336
rect 1903 11305 1915 11308
rect 1857 11299 1915 11305
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2682 11296 2688 11348
rect 2740 11336 2746 11348
rect 3418 11336 3424 11348
rect 2740 11308 3424 11336
rect 2740 11296 2746 11308
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 4982 11336 4988 11348
rect 4479 11308 4988 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 6181 11339 6239 11345
rect 6181 11305 6193 11339
rect 6227 11336 6239 11339
rect 7558 11336 7564 11348
rect 6227 11308 7564 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 1596 11240 2774 11268
rect 1596 11141 1624 11240
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 1719 11172 2329 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 2317 11169 2329 11172
rect 2363 11169 2375 11203
rect 2746 11200 2774 11240
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 6196 11268 6224 11299
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9306 11336 9312 11348
rect 9180 11308 9312 11336
rect 9180 11296 9186 11308
rect 9306 11296 9312 11308
rect 9364 11336 9370 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9364 11308 9689 11336
rect 9364 11296 9370 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 10594 11296 10600 11348
rect 10652 11296 10658 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 11514 11336 11520 11348
rect 10744 11308 11520 11336
rect 10744 11296 10750 11308
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11606 11296 11612 11348
rect 11664 11296 11670 11348
rect 11808 11308 13124 11336
rect 9490 11268 9496 11280
rect 3200 11240 6224 11268
rect 6380 11240 9496 11268
rect 3200 11228 3206 11240
rect 2746 11172 3280 11200
rect 2317 11163 2375 11169
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1581 11095 1639 11101
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2682 11132 2688 11144
rect 2455 11104 2688 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2240 11064 2268 11095
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 2792 11141 2820 11172
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 3142 11092 3148 11144
rect 3200 11092 3206 11144
rect 3252 11132 3280 11172
rect 3786 11160 3792 11212
rect 3844 11160 3850 11212
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4522 11200 4528 11212
rect 4111 11172 4528 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 6270 11160 6276 11212
rect 6328 11160 6334 11212
rect 3970 11132 3976 11144
rect 3252 11104 3976 11132
rect 3970 11092 3976 11104
rect 4028 11132 4034 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 4028 11104 4169 11132
rect 4028 11092 4034 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11132 4951 11135
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 4939 11104 6193 11132
rect 4939 11101 4951 11104
rect 4893 11095 4951 11101
rect 6181 11101 6193 11104
rect 6227 11132 6239 11135
rect 6380 11132 6408 11240
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11268 10563 11271
rect 10870 11268 10876 11280
rect 10551 11240 10876 11268
rect 10551 11237 10563 11240
rect 10505 11231 10563 11237
rect 10870 11228 10876 11240
rect 10928 11268 10934 11280
rect 11146 11268 11152 11280
rect 10928 11240 11152 11268
rect 10928 11228 10934 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 11808 11268 11836 11308
rect 11716 11240 11836 11268
rect 7024 11172 10640 11200
rect 6227 11104 6408 11132
rect 6457 11135 6515 11141
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6457 11101 6469 11135
rect 6503 11132 6515 11135
rect 6730 11132 6736 11144
rect 6503 11104 6736 11132
rect 6503 11101 6515 11104
rect 6457 11095 6515 11101
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7024 11141 7052 11172
rect 7009 11135 7067 11141
rect 7009 11101 7021 11135
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8904 11104 9137 11132
rect 8904 11092 8910 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2240 11036 2881 11064
rect 2869 11033 2881 11036
rect 2915 11033 2927 11067
rect 2869 11027 2927 11033
rect 2884 10996 2912 11027
rect 2958 11024 2964 11076
rect 3016 11073 3022 11076
rect 3016 11067 3065 11073
rect 3016 11033 3019 11067
rect 3053 11064 3065 11067
rect 3053 11036 3372 11064
rect 3053 11033 3065 11036
rect 3016 11027 3065 11033
rect 3016 11024 3022 11027
rect 3234 10996 3240 11008
rect 2884 10968 3240 10996
rect 3234 10956 3240 10968
rect 3292 10956 3298 11008
rect 3344 10996 3372 11036
rect 3418 11024 3424 11076
rect 3476 11024 3482 11076
rect 3605 11067 3663 11073
rect 3605 11033 3617 11067
rect 3651 11064 3663 11067
rect 4062 11064 4068 11076
rect 3651 11036 4068 11064
rect 3651 11033 3663 11036
rect 3605 11027 3663 11033
rect 3620 10996 3648 11027
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4246 11024 4252 11076
rect 4304 11073 4310 11076
rect 4304 11067 4332 11073
rect 4320 11033 4332 11067
rect 4304 11027 4332 11033
rect 4304 11024 4310 11027
rect 6270 11024 6276 11076
rect 6328 11064 6334 11076
rect 9217 11067 9275 11073
rect 9217 11064 9229 11067
rect 6328 11036 9229 11064
rect 6328 11024 6334 11036
rect 9217 11033 9229 11036
rect 9263 11064 9275 11067
rect 9674 11064 9680 11076
rect 9263 11036 9680 11064
rect 9263 11033 9275 11036
rect 9217 11027 9275 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 9784 11008 9812 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9916 11104 10425 11132
rect 9916 11092 9922 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10612 11132 10640 11172
rect 10686 11160 10692 11212
rect 10744 11160 10750 11212
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11716 11209 11744 11240
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11020 11172 11713 11200
rect 11020 11160 11026 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12250 11200 12256 11212
rect 11839 11172 12256 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12250 11160 12256 11172
rect 12308 11160 12314 11212
rect 12894 11200 12900 11212
rect 12406 11172 12900 11200
rect 10612 11104 11652 11132
rect 10413 11095 10471 11101
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 11517 11067 11575 11073
rect 11517 11064 11529 11067
rect 11388 11036 11529 11064
rect 11388 11024 11394 11036
rect 11517 11033 11529 11036
rect 11563 11033 11575 11067
rect 11624 11064 11652 11104
rect 11882 11092 11888 11144
rect 11940 11092 11946 11144
rect 12069 11135 12127 11141
rect 12069 11101 12081 11135
rect 12115 11132 12127 11135
rect 12406 11132 12434 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 12115 11104 12434 11132
rect 12115 11101 12127 11104
rect 12069 11095 12127 11101
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12710 11092 12716 11144
rect 12768 11092 12774 11144
rect 13096 11141 13124 11308
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 14902 11339 14960 11345
rect 14902 11336 14914 11339
rect 14792 11308 14914 11336
rect 14792 11296 14798 11308
rect 14902 11305 14914 11308
rect 14948 11305 14960 11339
rect 14902 11299 14960 11305
rect 15010 11296 15016 11348
rect 15068 11336 15074 11348
rect 16393 11339 16451 11345
rect 16393 11336 16405 11339
rect 15068 11308 16405 11336
rect 15068 11296 15074 11308
rect 16393 11305 16405 11308
rect 16439 11305 16451 11339
rect 16393 11299 16451 11305
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19576 11308 19717 11336
rect 19576 11296 19582 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 20530 11296 20536 11348
rect 20588 11336 20594 11348
rect 21545 11339 21603 11345
rect 21545 11336 21557 11339
rect 20588 11308 21557 11336
rect 20588 11296 20594 11308
rect 17218 11228 17224 11280
rect 17276 11268 17282 11280
rect 19613 11271 19671 11277
rect 17276 11240 17356 11268
rect 17276 11228 17282 11240
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 16482 11200 16488 11212
rect 13320 11172 16488 11200
rect 13320 11160 13326 11172
rect 16482 11160 16488 11172
rect 16540 11160 16546 11212
rect 17328 11200 17356 11240
rect 19613 11237 19625 11271
rect 19659 11268 19671 11271
rect 19797 11271 19855 11277
rect 19797 11268 19809 11271
rect 19659 11240 19809 11268
rect 19659 11237 19671 11240
rect 19613 11231 19671 11237
rect 19797 11237 19809 11240
rect 19843 11237 19855 11271
rect 20898 11268 20904 11280
rect 19797 11231 19855 11237
rect 20824 11240 20904 11268
rect 18785 11203 18843 11209
rect 18785 11200 18797 11203
rect 17328 11172 18797 11200
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11132 13139 11135
rect 13906 11132 13912 11144
rect 13127 11104 13912 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 12434 11064 12440 11076
rect 11624 11036 12440 11064
rect 11517 11027 11575 11033
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 13004 11064 13032 11095
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 14274 11092 14280 11144
rect 14332 11132 14338 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14332 11104 14657 11132
rect 14332 11092 14338 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 16666 11092 16672 11144
rect 16724 11092 16730 11144
rect 17034 11092 17040 11144
rect 17092 11092 17098 11144
rect 17328 11141 17356 11172
rect 18785 11169 18797 11172
rect 18831 11169 18843 11203
rect 18785 11163 18843 11169
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11101 17371 11135
rect 17313 11095 17371 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 13004 11036 13124 11064
rect 16146 11036 16589 11064
rect 13096 11008 13124 11036
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 17236 11064 17264 11095
rect 17512 11064 17540 11095
rect 17586 11092 17592 11144
rect 17644 11092 17650 11144
rect 17773 11135 17831 11141
rect 17773 11101 17785 11135
rect 17819 11132 17831 11135
rect 17862 11132 17868 11144
rect 17819 11104 17868 11132
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18564 11104 18705 11132
rect 18564 11092 18570 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 18693 11095 18751 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 19058 11132 19064 11144
rect 18923 11104 19064 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 17681 11067 17739 11073
rect 17681 11064 17693 11067
rect 17236 11036 17693 11064
rect 16577 11027 16635 11033
rect 17681 11033 17693 11036
rect 17727 11033 17739 11067
rect 18708 11064 18736 11095
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20257 11135 20315 11141
rect 20257 11101 20269 11135
rect 20303 11132 20315 11135
rect 20303 11104 20337 11132
rect 20303 11101 20315 11104
rect 20257 11095 20315 11101
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18708 11036 19257 11064
rect 17681 11027 17739 11033
rect 19245 11033 19257 11036
rect 19291 11033 19303 11067
rect 19245 11027 19303 11033
rect 19794 11024 19800 11076
rect 19852 11064 19858 11076
rect 20272 11064 20300 11095
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 20622 11092 20628 11144
rect 20680 11092 20686 11144
rect 20824 11141 20852 11240
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 21008 11141 21036 11308
rect 21545 11305 21557 11308
rect 21591 11305 21603 11339
rect 21545 11299 21603 11305
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 22833 11339 22891 11345
rect 22833 11336 22845 11339
rect 22612 11308 22845 11336
rect 22612 11296 22618 11308
rect 22833 11305 22845 11308
rect 22879 11305 22891 11339
rect 22833 11299 22891 11305
rect 23014 11296 23020 11348
rect 23072 11296 23078 11348
rect 27522 11296 27528 11348
rect 27580 11336 27586 11348
rect 28077 11339 28135 11345
rect 28077 11336 28089 11339
rect 27580 11308 28089 11336
rect 27580 11296 27586 11308
rect 28077 11305 28089 11308
rect 28123 11305 28135 11339
rect 28077 11299 28135 11305
rect 28813 11339 28871 11345
rect 28813 11305 28825 11339
rect 28859 11336 28871 11339
rect 28994 11336 29000 11348
rect 28859 11308 29000 11336
rect 28859 11305 28871 11308
rect 28813 11299 28871 11305
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 21269 11271 21327 11277
rect 21269 11237 21281 11271
rect 21315 11268 21327 11271
rect 21726 11268 21732 11280
rect 21315 11240 21732 11268
rect 21315 11237 21327 11240
rect 21269 11231 21327 11237
rect 21726 11228 21732 11240
rect 21784 11228 21790 11280
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 21968 11240 25636 11268
rect 21968 11228 21974 11240
rect 22005 11203 22063 11209
rect 22005 11169 22017 11203
rect 22051 11200 22063 11203
rect 22278 11200 22284 11212
rect 22051 11172 22284 11200
rect 22051 11169 22063 11172
rect 22005 11163 22063 11169
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 22462 11160 22468 11212
rect 22520 11200 22526 11212
rect 22741 11203 22799 11209
rect 22741 11200 22753 11203
rect 22520 11172 22753 11200
rect 22520 11160 22526 11172
rect 22741 11169 22753 11172
rect 22787 11169 22799 11203
rect 22741 11163 22799 11169
rect 22830 11160 22836 11212
rect 22888 11200 22894 11212
rect 23201 11203 23259 11209
rect 22888 11172 23152 11200
rect 22888 11160 22894 11172
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11101 20867 11135
rect 20809 11095 20867 11101
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11101 20959 11135
rect 20901 11095 20959 11101
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11101 21051 11135
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20993 11095 21051 11101
rect 21284 11104 21373 11132
rect 20349 11067 20407 11073
rect 20349 11064 20361 11067
rect 19852 11036 20361 11064
rect 19852 11024 19858 11036
rect 20349 11033 20361 11036
rect 20395 11033 20407 11067
rect 20640 11064 20668 11092
rect 20916 11064 20944 11095
rect 21284 11076 21312 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21542 11092 21548 11144
rect 21600 11092 21606 11144
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 21744 11104 22109 11132
rect 21266 11064 21272 11076
rect 20640 11036 20852 11064
rect 20916 11036 21272 11064
rect 20349 11027 20407 11033
rect 3344 10968 3648 10996
rect 6638 10956 6644 11008
rect 6696 10956 6702 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7374 10996 7380 11008
rect 7156 10968 7380 10996
rect 7156 10956 7162 10968
rect 7374 10956 7380 10968
rect 7432 10996 7438 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 7432 10968 8309 10996
rect 7432 10956 7438 10968
rect 8297 10965 8309 10968
rect 8343 10965 8355 10999
rect 8297 10959 8355 10965
rect 8941 10999 8999 11005
rect 8941 10965 8953 10999
rect 8987 10996 8999 10999
rect 9122 10996 9128 11008
rect 8987 10968 9128 10996
rect 8987 10965 8999 10968
rect 8941 10959 8999 10965
rect 9122 10956 9128 10968
rect 9180 10956 9186 11008
rect 9766 10956 9772 11008
rect 9824 10996 9830 11008
rect 11698 10996 11704 11008
rect 9824 10968 11704 10996
rect 9824 10956 9830 10968
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12897 10999 12955 11005
rect 12897 10996 12909 10999
rect 12584 10968 12909 10996
rect 12584 10956 12590 10968
rect 12897 10965 12909 10968
rect 12943 10996 12955 10999
rect 12986 10996 12992 11008
rect 12943 10968 12992 10996
rect 12943 10965 12955 10968
rect 12897 10959 12955 10965
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 13173 10999 13231 11005
rect 13173 10996 13185 10999
rect 13136 10968 13185 10996
rect 13136 10956 13142 10968
rect 13173 10965 13185 10968
rect 13219 10965 13231 10999
rect 13173 10959 13231 10965
rect 17129 10999 17187 11005
rect 17129 10965 17141 10999
rect 17175 10996 17187 10999
rect 17310 10996 17316 11008
rect 17175 10968 17316 10996
rect 17175 10965 17187 10968
rect 17129 10959 17187 10965
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 17402 10956 17408 11008
rect 17460 10956 17466 11008
rect 20162 10956 20168 11008
rect 20220 10956 20226 11008
rect 20824 10996 20852 11036
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21634 11024 21640 11076
rect 21692 11024 21698 11076
rect 21085 10999 21143 11005
rect 21085 10996 21097 10999
rect 20824 10968 21097 10996
rect 21085 10965 21097 10968
rect 21131 10996 21143 10999
rect 21744 10996 21772 11104
rect 22097 11101 22109 11104
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 22373 11135 22431 11141
rect 22373 11101 22385 11135
rect 22419 11132 22431 11135
rect 22848 11132 22876 11160
rect 22419 11104 22876 11132
rect 23017 11135 23075 11141
rect 22419 11101 22431 11104
rect 22373 11095 22431 11101
rect 23017 11101 23029 11135
rect 23063 11101 23075 11135
rect 23124 11132 23152 11172
rect 23201 11169 23213 11203
rect 23247 11200 23259 11203
rect 23474 11200 23480 11212
rect 23247 11172 23480 11200
rect 23247 11169 23259 11172
rect 23201 11163 23259 11169
rect 23474 11160 23480 11172
rect 23532 11200 23538 11212
rect 24486 11200 24492 11212
rect 23532 11172 24492 11200
rect 23532 11160 23538 11172
rect 24486 11160 24492 11172
rect 24544 11160 24550 11212
rect 25608 11200 25636 11240
rect 27982 11228 27988 11280
rect 28040 11228 28046 11280
rect 29181 11271 29239 11277
rect 29181 11237 29193 11271
rect 29227 11237 29239 11271
rect 29181 11231 29239 11237
rect 29196 11200 29224 11231
rect 25608 11172 29224 11200
rect 23293 11135 23351 11141
rect 23293 11132 23305 11135
rect 23124 11104 23305 11132
rect 23017 11095 23075 11101
rect 23293 11101 23305 11104
rect 23339 11101 23351 11135
rect 23293 11095 23351 11101
rect 26053 11135 26111 11141
rect 26053 11101 26065 11135
rect 26099 11132 26111 11135
rect 26142 11132 26148 11144
rect 26099 11104 26148 11132
rect 26099 11101 26111 11104
rect 26053 11095 26111 11101
rect 21818 11024 21824 11076
rect 21876 11024 21882 11076
rect 23032 11064 23060 11095
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 26329 11135 26387 11141
rect 26329 11101 26341 11135
rect 26375 11132 26387 11135
rect 26418 11132 26424 11144
rect 26375 11104 26424 11132
rect 26375 11101 26387 11104
rect 26329 11095 26387 11101
rect 26418 11092 26424 11104
rect 26476 11092 26482 11144
rect 27617 11135 27675 11141
rect 27617 11101 27629 11135
rect 27663 11132 27675 11135
rect 27798 11132 27804 11144
rect 27663 11104 27804 11132
rect 27663 11101 27675 11104
rect 27617 11095 27675 11101
rect 27798 11092 27804 11104
rect 27856 11092 27862 11144
rect 28074 11092 28080 11144
rect 28132 11092 28138 11144
rect 28258 11092 28264 11144
rect 28316 11092 28322 11144
rect 28902 11092 28908 11144
rect 28960 11092 28966 11144
rect 29362 11092 29368 11144
rect 29420 11092 29426 11144
rect 23198 11064 23204 11076
rect 23032 11036 23204 11064
rect 23198 11024 23204 11036
rect 23256 11024 23262 11076
rect 26237 11067 26295 11073
rect 26237 11033 26249 11067
rect 26283 11033 26295 11067
rect 26237 11027 26295 11033
rect 21131 10968 21772 10996
rect 21131 10965 21143 10968
rect 21085 10959 21143 10965
rect 25314 10956 25320 11008
rect 25372 10996 25378 11008
rect 25961 10999 26019 11005
rect 25961 10996 25973 10999
rect 25372 10968 25973 10996
rect 25372 10956 25378 10968
rect 25961 10965 25973 10968
rect 26007 10965 26019 10999
rect 26252 10996 26280 11027
rect 27430 11024 27436 11076
rect 27488 11024 27494 11076
rect 27709 11067 27767 11073
rect 27709 11033 27721 11067
rect 27755 11064 27767 11067
rect 28276 11064 28304 11092
rect 27755 11036 28304 11064
rect 27755 11033 27767 11036
rect 27709 11027 27767 11033
rect 26326 10996 26332 11008
rect 26252 10968 26332 10996
rect 25961 10959 26019 10965
rect 26326 10956 26332 10968
rect 26384 10956 26390 11008
rect 27798 10956 27804 11008
rect 27856 10956 27862 11008
rect 1104 10906 29716 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 29716 10906
rect 1104 10832 29716 10854
rect 3513 10795 3571 10801
rect 3513 10761 3525 10795
rect 3559 10792 3571 10795
rect 4246 10792 4252 10804
rect 3559 10764 4252 10792
rect 3559 10761 3571 10764
rect 3513 10755 3571 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 7101 10795 7159 10801
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7190 10792 7196 10804
rect 7147 10764 7196 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7800 10764 8125 10792
rect 7800 10752 7806 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 8938 10752 8944 10804
rect 8996 10792 9002 10804
rect 9766 10792 9772 10804
rect 8996 10764 9772 10792
rect 8996 10752 9002 10764
rect 9766 10752 9772 10764
rect 9824 10752 9830 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 12952 10764 13768 10792
rect 12952 10752 12958 10764
rect 842 10684 848 10736
rect 900 10724 906 10736
rect 1489 10727 1547 10733
rect 1489 10724 1501 10727
rect 900 10696 1501 10724
rect 900 10684 906 10696
rect 1489 10693 1501 10696
rect 1535 10693 1547 10727
rect 1489 10687 1547 10693
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 3605 10727 3663 10733
rect 3605 10724 3617 10727
rect 2740 10696 3617 10724
rect 2740 10684 2746 10696
rect 3605 10693 3617 10696
rect 3651 10693 3663 10727
rect 3605 10687 3663 10693
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 6696 10696 6745 10724
rect 6696 10684 6702 10696
rect 6733 10693 6745 10696
rect 6779 10693 6791 10727
rect 8846 10724 8852 10736
rect 6733 10687 6791 10693
rect 8404 10696 8852 10724
rect 1670 10616 1676 10668
rect 1728 10616 1734 10668
rect 2590 10616 2596 10668
rect 2648 10616 2654 10668
rect 2777 10659 2835 10665
rect 2777 10625 2789 10659
rect 2823 10656 2835 10659
rect 2866 10656 2872 10668
rect 2823 10628 2872 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3053 10659 3111 10665
rect 3053 10656 3065 10659
rect 3007 10628 3065 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3053 10625 3065 10628
rect 3099 10656 3111 10659
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3099 10628 3801 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3970 10616 3976 10668
rect 4028 10616 4034 10668
rect 4522 10616 4528 10668
rect 4580 10656 4586 10668
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4580 10628 5089 10656
rect 4580 10616 4586 10628
rect 5077 10625 5089 10628
rect 5123 10656 5135 10659
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5123 10628 5457 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6604 10628 6929 10656
rect 6604 10616 6610 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 8404 10665 8432 10696
rect 8846 10684 8852 10696
rect 8904 10684 8910 10736
rect 10597 10727 10655 10733
rect 9692 10696 10548 10724
rect 9692 10668 9720 10696
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7156 10628 7389 10656
rect 7156 10616 7162 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5718 10588 5724 10600
rect 5399 10560 5724 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 8680 10588 8708 10619
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 9180 10628 9229 10656
rect 9180 10616 9186 10628
rect 9217 10625 9229 10628
rect 9263 10625 9275 10659
rect 9217 10619 9275 10625
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9398 10616 9404 10668
rect 9456 10616 9462 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 9674 10656 9680 10668
rect 9631 10628 9680 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10625 10471 10659
rect 10520 10656 10548 10696
rect 10597 10693 10609 10727
rect 10643 10724 10655 10727
rect 11330 10724 11336 10736
rect 10643 10696 11336 10724
rect 10643 10693 10655 10696
rect 10597 10687 10655 10693
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 12434 10684 12440 10736
rect 12492 10724 12498 10736
rect 13262 10724 13268 10736
rect 12492 10696 13268 10724
rect 12492 10684 12498 10696
rect 13262 10684 13268 10696
rect 13320 10684 13326 10736
rect 13354 10684 13360 10736
rect 13412 10684 13418 10736
rect 10689 10659 10747 10665
rect 10689 10656 10701 10659
rect 10520 10628 10701 10656
rect 10413 10619 10471 10625
rect 10689 10625 10701 10628
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 10870 10656 10876 10668
rect 10827 10628 10876 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 9140 10588 9168 10616
rect 8680 10560 9168 10588
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 10428 10588 10456 10619
rect 10594 10588 10600 10600
rect 9548 10560 10600 10588
rect 9548 10548 9554 10560
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10704 10588 10732 10619
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 13136 10628 13553 10656
rect 13136 10616 13142 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13630 10616 13636 10668
rect 13688 10616 13694 10668
rect 13740 10665 13768 10764
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14642 10792 14648 10804
rect 14148 10764 14648 10792
rect 14148 10752 14154 10764
rect 14642 10752 14648 10764
rect 14700 10752 14706 10804
rect 18877 10795 18935 10801
rect 18877 10761 18889 10795
rect 18923 10792 18935 10795
rect 19058 10792 19064 10804
rect 18923 10764 19064 10792
rect 18923 10761 18935 10764
rect 18877 10755 18935 10761
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19153 10795 19211 10801
rect 19153 10761 19165 10795
rect 19199 10792 19211 10795
rect 19242 10792 19248 10804
rect 19199 10764 19248 10792
rect 19199 10761 19211 10764
rect 19153 10755 19211 10761
rect 19242 10752 19248 10764
rect 19300 10752 19306 10804
rect 19689 10795 19747 10801
rect 19689 10761 19701 10795
rect 19735 10792 19747 10795
rect 19794 10792 19800 10804
rect 19735 10764 19800 10792
rect 19735 10761 19747 10764
rect 19689 10755 19747 10761
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 20073 10795 20131 10801
rect 20073 10761 20085 10795
rect 20119 10792 20131 10795
rect 20162 10792 20168 10804
rect 20119 10764 20168 10792
rect 20119 10761 20131 10764
rect 20073 10755 20131 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21266 10792 21272 10804
rect 21131 10764 21272 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21266 10752 21272 10764
rect 21324 10752 21330 10804
rect 21542 10752 21548 10804
rect 21600 10792 21606 10804
rect 21913 10795 21971 10801
rect 21913 10792 21925 10795
rect 21600 10764 21925 10792
rect 21600 10752 21606 10764
rect 21913 10761 21925 10764
rect 21959 10761 21971 10795
rect 21913 10755 21971 10761
rect 26234 10752 26240 10804
rect 26292 10792 26298 10804
rect 26789 10795 26847 10801
rect 26789 10792 26801 10795
rect 26292 10764 26801 10792
rect 26292 10752 26298 10764
rect 26789 10761 26801 10764
rect 26835 10792 26847 10795
rect 27430 10792 27436 10804
rect 26835 10764 27436 10792
rect 26835 10761 26847 10764
rect 26789 10755 26847 10761
rect 27430 10752 27436 10764
rect 27488 10792 27494 10804
rect 27488 10764 27568 10792
rect 27488 10752 27494 10764
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 14918 10724 14924 10736
rect 13964 10696 14924 10724
rect 13964 10684 13970 10696
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 17954 10724 17960 10736
rect 16960 10696 17960 10724
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13771 10628 14013 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 14001 10625 14013 10628
rect 14047 10656 14059 10659
rect 15010 10656 15016 10668
rect 14047 10628 15016 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 16960 10665 16988 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18414 10684 18420 10736
rect 18472 10724 18478 10736
rect 19889 10727 19947 10733
rect 18472 10696 19840 10724
rect 18472 10684 18478 10696
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 10962 10588 10968 10600
rect 10704 10560 10968 10588
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 16853 10591 16911 10597
rect 12406 10560 16804 10588
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 3329 10523 3387 10529
rect 3329 10520 3341 10523
rect 3292 10492 3341 10520
rect 3292 10480 3298 10492
rect 3329 10489 3341 10492
rect 3375 10489 3387 10523
rect 3329 10483 3387 10489
rect 5261 10523 5319 10529
rect 5261 10489 5273 10523
rect 5307 10520 5319 10523
rect 5537 10523 5595 10529
rect 5537 10520 5549 10523
rect 5307 10492 5549 10520
rect 5307 10489 5319 10492
rect 5261 10483 5319 10489
rect 5368 10464 5396 10492
rect 5537 10489 5549 10492
rect 5583 10489 5595 10523
rect 5537 10483 5595 10489
rect 7190 10480 7196 10532
rect 7248 10520 7254 10532
rect 12406 10520 12434 10560
rect 7248 10492 12434 10520
rect 16776 10520 16804 10560
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 17034 10588 17040 10600
rect 16899 10560 17040 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 17034 10548 17040 10560
rect 17092 10588 17098 10600
rect 17236 10588 17264 10619
rect 17402 10616 17408 10668
rect 17460 10616 17466 10668
rect 17862 10616 17868 10668
rect 17920 10616 17926 10668
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 17092 10560 17264 10588
rect 18800 10588 18828 10619
rect 18874 10616 18880 10668
rect 18932 10662 18938 10668
rect 19076 10665 19104 10696
rect 18969 10662 19027 10665
rect 18932 10659 19027 10662
rect 18932 10634 18981 10659
rect 18932 10616 18938 10634
rect 18969 10625 18981 10634
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19245 10659 19303 10665
rect 19245 10625 19257 10659
rect 19291 10656 19303 10659
rect 19702 10656 19708 10668
rect 19291 10628 19708 10656
rect 19291 10625 19303 10628
rect 19245 10619 19303 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19812 10656 19840 10696
rect 19889 10693 19901 10727
rect 19935 10724 19947 10727
rect 19978 10724 19984 10736
rect 19935 10696 19984 10724
rect 19935 10693 19947 10696
rect 19889 10687 19947 10693
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 20441 10727 20499 10733
rect 20441 10724 20453 10727
rect 20088 10696 20453 10724
rect 20088 10656 20116 10696
rect 20441 10693 20453 10696
rect 20487 10693 20499 10727
rect 20441 10687 20499 10693
rect 19812 10628 20116 10656
rect 20254 10616 20260 10668
rect 20312 10616 20318 10668
rect 20456 10656 20484 10687
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 20772 10696 22876 10724
rect 20772 10684 20778 10696
rect 21174 10656 21180 10668
rect 20456 10628 21180 10656
rect 21174 10616 21180 10628
rect 21232 10656 21238 10668
rect 21269 10659 21327 10665
rect 21269 10656 21281 10659
rect 21232 10628 21281 10656
rect 21232 10616 21238 10628
rect 21269 10625 21281 10628
rect 21315 10656 21327 10659
rect 21634 10656 21640 10668
rect 21315 10628 21640 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 21634 10616 21640 10628
rect 21692 10656 21698 10668
rect 22848 10665 22876 10696
rect 24118 10684 24124 10736
rect 24176 10684 24182 10736
rect 25314 10684 25320 10736
rect 25372 10684 25378 10736
rect 26326 10684 26332 10736
rect 26384 10684 26390 10736
rect 27540 10733 27568 10764
rect 27798 10733 27804 10736
rect 27525 10727 27583 10733
rect 27525 10693 27537 10727
rect 27571 10693 27583 10727
rect 27525 10687 27583 10693
rect 27741 10727 27804 10733
rect 27741 10693 27753 10727
rect 27787 10693 27804 10727
rect 27741 10687 27804 10693
rect 27798 10684 27804 10687
rect 27856 10684 27862 10736
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21692 10628 21833 10656
rect 21692 10616 21698 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 22005 10659 22063 10665
rect 22005 10625 22017 10659
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 20070 10588 20076 10600
rect 18800 10560 20076 10588
rect 17092 10548 17098 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 21453 10591 21511 10597
rect 21453 10557 21465 10591
rect 21499 10588 21511 10591
rect 22020 10588 22048 10619
rect 27890 10616 27896 10668
rect 27948 10656 27954 10668
rect 27985 10659 28043 10665
rect 27985 10656 27997 10659
rect 27948 10628 27997 10656
rect 27948 10616 27954 10628
rect 27985 10625 27997 10628
rect 28031 10625 28043 10659
rect 27985 10619 28043 10625
rect 28169 10659 28227 10665
rect 28169 10625 28181 10659
rect 28215 10625 28227 10659
rect 28169 10619 28227 10625
rect 22370 10588 22376 10600
rect 21499 10560 22376 10588
rect 21499 10557 21511 10560
rect 21453 10551 21511 10557
rect 22370 10548 22376 10560
rect 22428 10548 22434 10600
rect 23106 10548 23112 10600
rect 23164 10548 23170 10600
rect 23198 10548 23204 10600
rect 23256 10588 23262 10600
rect 24857 10591 24915 10597
rect 24857 10588 24869 10591
rect 23256 10560 24869 10588
rect 23256 10548 23262 10560
rect 24857 10557 24869 10560
rect 24903 10557 24915 10591
rect 24857 10551 24915 10557
rect 25038 10548 25044 10600
rect 25096 10548 25102 10600
rect 28074 10588 28080 10600
rect 27908 10560 28080 10588
rect 18138 10520 18144 10532
rect 16776 10492 18144 10520
rect 7248 10480 7254 10492
rect 18138 10480 18144 10492
rect 18196 10480 18202 10532
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 19521 10523 19579 10529
rect 19521 10520 19533 10523
rect 18564 10492 19533 10520
rect 18564 10480 18570 10492
rect 19521 10489 19533 10492
rect 19567 10489 19579 10523
rect 21542 10520 21548 10532
rect 19521 10483 19579 10489
rect 19628 10492 21548 10520
rect 4890 10412 4896 10464
rect 4948 10412 4954 10464
rect 5350 10412 5356 10464
rect 5408 10412 5414 10464
rect 5442 10412 5448 10464
rect 5500 10412 5506 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8297 10455 8355 10461
rect 8297 10452 8309 10455
rect 7984 10424 8309 10452
rect 7984 10412 7990 10424
rect 8297 10421 8309 10424
rect 8343 10421 8355 10455
rect 8297 10415 8355 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9306 10452 9312 10464
rect 8904 10424 9312 10452
rect 8904 10412 8910 10424
rect 9306 10412 9312 10424
rect 9364 10452 9370 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9364 10424 9413 10452
rect 9364 10412 9370 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10686 10452 10692 10464
rect 10284 10424 10692 10452
rect 10284 10412 10290 10424
rect 10686 10412 10692 10424
rect 10744 10452 10750 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10744 10424 10977 10452
rect 10744 10412 10750 10424
rect 10965 10421 10977 10424
rect 11011 10421 11023 10455
rect 10965 10415 11023 10421
rect 11790 10412 11796 10464
rect 11848 10412 11854 10464
rect 12250 10412 12256 10464
rect 12308 10452 12314 10464
rect 13814 10452 13820 10464
rect 12308 10424 13820 10452
rect 12308 10412 12314 10424
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 17402 10412 17408 10464
rect 17460 10412 17466 10464
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 19426 10452 19432 10464
rect 18932 10424 19432 10452
rect 18932 10412 18938 10424
rect 19426 10412 19432 10424
rect 19484 10452 19490 10464
rect 19628 10452 19656 10492
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 27908 10529 27936 10560
rect 28074 10548 28080 10560
rect 28132 10588 28138 10600
rect 28184 10588 28212 10619
rect 28132 10560 28212 10588
rect 28132 10548 28138 10560
rect 27893 10523 27951 10529
rect 27893 10489 27905 10523
rect 27939 10489 27951 10523
rect 27893 10483 27951 10489
rect 19484 10424 19656 10452
rect 19705 10455 19763 10461
rect 19484 10412 19490 10424
rect 19705 10421 19717 10455
rect 19751 10452 19763 10455
rect 20162 10452 20168 10464
rect 19751 10424 20168 10452
rect 19751 10421 19763 10424
rect 19705 10415 19763 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 27706 10412 27712 10464
rect 27764 10412 27770 10464
rect 27982 10412 27988 10464
rect 28040 10412 28046 10464
rect 1104 10362 29716 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 29716 10362
rect 1104 10288 29716 10310
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4157 10251 4215 10257
rect 4157 10248 4169 10251
rect 4028 10220 4169 10248
rect 4028 10208 4034 10220
rect 4157 10217 4169 10220
rect 4203 10217 4215 10251
rect 4157 10211 4215 10217
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 6365 10251 6423 10257
rect 6365 10248 6377 10251
rect 5776 10220 6377 10248
rect 5776 10208 5782 10220
rect 6365 10217 6377 10220
rect 6411 10217 6423 10251
rect 6365 10211 6423 10217
rect 7006 10208 7012 10260
rect 7064 10208 7070 10260
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 10502 10248 10508 10260
rect 9723 10220 10508 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10781 10251 10839 10257
rect 10781 10217 10793 10251
rect 10827 10248 10839 10251
rect 10870 10248 10876 10260
rect 10827 10220 10876 10248
rect 10827 10217 10839 10220
rect 10781 10211 10839 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12802 10208 12808 10260
rect 12860 10208 12866 10260
rect 13722 10208 13728 10260
rect 13780 10208 13786 10260
rect 13909 10251 13967 10257
rect 13909 10217 13921 10251
rect 13955 10248 13967 10251
rect 15669 10251 15727 10257
rect 15669 10248 15681 10251
rect 13955 10220 15681 10248
rect 13955 10217 13967 10220
rect 13909 10211 13967 10217
rect 15669 10217 15681 10220
rect 15715 10217 15727 10251
rect 15669 10211 15727 10217
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 17034 10248 17040 10260
rect 16623 10220 17040 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 17034 10208 17040 10220
rect 17092 10248 17098 10260
rect 17497 10251 17555 10257
rect 17497 10248 17509 10251
rect 17092 10220 17509 10248
rect 17092 10208 17098 10220
rect 17497 10217 17509 10220
rect 17543 10217 17555 10251
rect 17497 10211 17555 10217
rect 18138 10208 18144 10260
rect 18196 10208 18202 10260
rect 18322 10208 18328 10260
rect 18380 10248 18386 10260
rect 19334 10248 19340 10260
rect 18380 10220 18920 10248
rect 18380 10208 18386 10220
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 6825 10183 6883 10189
rect 6825 10180 6837 10183
rect 5408 10152 6837 10180
rect 5408 10140 5414 10152
rect 6825 10149 6837 10152
rect 6871 10149 6883 10183
rect 6825 10143 6883 10149
rect 12713 10183 12771 10189
rect 12713 10149 12725 10183
rect 12759 10180 12771 10183
rect 12894 10180 12900 10192
rect 12759 10152 12900 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13262 10140 13268 10192
rect 13320 10180 13326 10192
rect 13630 10180 13636 10192
rect 13320 10152 13636 10180
rect 13320 10140 13326 10152
rect 13630 10140 13636 10152
rect 13688 10180 13694 10192
rect 14185 10183 14243 10189
rect 14185 10180 14197 10183
rect 13688 10152 14197 10180
rect 13688 10140 13694 10152
rect 14185 10149 14197 10152
rect 14231 10149 14243 10183
rect 14185 10143 14243 10149
rect 17681 10183 17739 10189
rect 17681 10149 17693 10183
rect 17727 10149 17739 10183
rect 17681 10143 17739 10149
rect 4798 10112 4804 10124
rect 4632 10084 4804 10112
rect 4632 10053 4660 10084
rect 4798 10072 4804 10084
rect 4856 10112 4862 10124
rect 6362 10112 6368 10124
rect 4856 10084 6368 10112
rect 4856 10072 4862 10084
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6420 10084 6745 10112
rect 6420 10072 6426 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 14274 10112 14280 10124
rect 6733 10075 6791 10081
rect 12406 10084 14280 10112
rect 4341 10047 4399 10053
rect 4341 10013 4353 10047
rect 4387 10013 4399 10047
rect 4341 10007 4399 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 4356 9976 4384 10007
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5442 10044 5448 10056
rect 5123 10016 5448 10044
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8754 10044 8760 10056
rect 8067 10016 8760 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 9950 10004 9956 10056
rect 10008 10004 10014 10056
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 10100 10016 10149 10044
rect 10100 10004 10106 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 4908 9976 4936 10004
rect 4356 9948 4936 9976
rect 7190 9936 7196 9988
rect 7248 9936 7254 9988
rect 10520 9976 10548 10007
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10873 10047 10931 10053
rect 10873 10013 10885 10047
rect 10919 10044 10931 10047
rect 10962 10044 10968 10056
rect 10919 10016 10968 10044
rect 10919 10013 10931 10016
rect 10873 10007 10931 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11790 10004 11796 10056
rect 11848 10044 11854 10056
rect 12406 10044 12434 10084
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 14332 10084 15945 10112
rect 14332 10072 14338 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 17494 10112 17500 10124
rect 16347 10084 17500 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 17696 10112 17724 10143
rect 17862 10140 17868 10192
rect 17920 10180 17926 10192
rect 18892 10180 18920 10220
rect 19306 10208 19340 10248
rect 19392 10208 19398 10260
rect 19521 10251 19579 10257
rect 19521 10217 19533 10251
rect 19567 10217 19579 10251
rect 19521 10211 19579 10217
rect 19306 10180 19334 10208
rect 17920 10152 18828 10180
rect 18892 10152 19334 10180
rect 17920 10140 17926 10152
rect 18800 10112 18828 10152
rect 19337 10115 19395 10121
rect 19337 10112 19349 10115
rect 17696 10084 18736 10112
rect 18800 10084 19349 10112
rect 11848 10016 12434 10044
rect 11848 10004 11854 10016
rect 12618 10004 12624 10056
rect 12676 10044 12682 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12676 10016 12817 10044
rect 12676 10004 12682 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 16206 10004 16212 10056
rect 16264 10044 16270 10056
rect 16264 10016 18092 10044
rect 16264 10004 16270 10016
rect 11330 9976 11336 9988
rect 10520 9948 11336 9976
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 12529 9979 12587 9985
rect 12529 9976 12541 9979
rect 11664 9948 12541 9976
rect 11664 9936 11670 9948
rect 12529 9945 12541 9948
rect 12575 9945 12587 9979
rect 12529 9939 12587 9945
rect 13078 9936 13084 9988
rect 13136 9936 13142 9988
rect 13541 9979 13599 9985
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13998 9976 14004 9988
rect 13587 9948 14004 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 13998 9936 14004 9948
rect 14056 9976 14062 9988
rect 14366 9976 14372 9988
rect 14056 9948 14372 9976
rect 14056 9936 14062 9948
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 14918 9936 14924 9988
rect 14976 9936 14982 9988
rect 17310 9936 17316 9988
rect 17368 9936 17374 9988
rect 4522 9868 4528 9920
rect 4580 9868 4586 9920
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 4985 9911 5043 9917
rect 4985 9908 4997 9911
rect 4856 9880 4997 9908
rect 4856 9868 4862 9880
rect 4985 9877 4997 9880
rect 5031 9877 5043 9911
rect 4985 9871 5043 9877
rect 6993 9911 7051 9917
rect 6993 9877 7005 9911
rect 7039 9908 7051 9911
rect 7282 9908 7288 9920
rect 7039 9880 7288 9908
rect 7039 9877 7051 9880
rect 6993 9871 7051 9877
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 10321 9911 10379 9917
rect 10321 9908 10333 9911
rect 10192 9880 10333 9908
rect 10192 9868 10198 9880
rect 10321 9877 10333 9880
rect 10367 9877 10379 9911
rect 10321 9871 10379 9877
rect 13449 9911 13507 9917
rect 13449 9877 13461 9911
rect 13495 9908 13507 9911
rect 13741 9911 13799 9917
rect 13741 9908 13753 9911
rect 13495 9880 13753 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13741 9877 13753 9880
rect 13787 9877 13799 9911
rect 13741 9871 13799 9877
rect 17523 9911 17581 9917
rect 17523 9877 17535 9911
rect 17569 9908 17581 9911
rect 17862 9908 17868 9920
rect 17569 9880 17868 9908
rect 17569 9877 17581 9880
rect 17523 9871 17581 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18064 9908 18092 10016
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 18708 10053 18736 10084
rect 19337 10081 19349 10084
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19536 10112 19564 10211
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19668 10220 19717 10248
rect 19668 10208 19674 10220
rect 19705 10217 19717 10220
rect 19751 10248 19763 10251
rect 19886 10248 19892 10260
rect 19751 10220 19892 10248
rect 19751 10217 19763 10220
rect 19705 10211 19763 10217
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 22833 10251 22891 10257
rect 22833 10217 22845 10251
rect 22879 10248 22891 10251
rect 23106 10248 23112 10260
rect 22879 10220 23112 10248
rect 22879 10217 22891 10220
rect 22833 10211 22891 10217
rect 23106 10208 23112 10220
rect 23164 10208 23170 10260
rect 24118 10208 24124 10260
rect 24176 10208 24182 10260
rect 26418 10248 26424 10260
rect 24228 10220 26424 10248
rect 19484 10084 19564 10112
rect 19484 10072 19490 10084
rect 21634 10072 21640 10124
rect 21692 10072 21698 10124
rect 23198 10072 23204 10124
rect 23256 10112 23262 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 23256 10084 23305 10112
rect 23256 10072 23262 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23477 10115 23535 10121
rect 23477 10081 23489 10115
rect 23523 10112 23535 10115
rect 23658 10112 23664 10124
rect 23523 10084 23664 10112
rect 23523 10081 23535 10084
rect 23477 10075 23535 10081
rect 23658 10072 23664 10084
rect 23716 10072 23722 10124
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10013 18751 10047
rect 19521 10047 19579 10053
rect 19521 10044 19533 10047
rect 18693 10007 18751 10013
rect 18800 10016 19533 10044
rect 18414 9936 18420 9988
rect 18472 9936 18478 9988
rect 18800 9908 18828 10016
rect 19521 10013 19533 10016
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 19981 10047 20039 10053
rect 19981 10044 19993 10047
rect 19760 10016 19993 10044
rect 19760 10004 19766 10016
rect 19981 10013 19993 10016
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 21726 10004 21732 10056
rect 21784 10004 21790 10056
rect 24228 10053 24256 10220
rect 26418 10208 26424 10220
rect 26476 10208 26482 10260
rect 27525 10251 27583 10257
rect 27525 10217 27537 10251
rect 27571 10248 27583 10251
rect 27890 10248 27896 10260
rect 27571 10220 27896 10248
rect 27571 10217 27583 10220
rect 27525 10211 27583 10217
rect 27890 10208 27896 10220
rect 27948 10208 27954 10260
rect 26068 10152 27292 10180
rect 26068 10121 26096 10152
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10081 26111 10115
rect 26053 10075 26111 10081
rect 26326 10072 26332 10124
rect 26384 10072 26390 10124
rect 24213 10047 24271 10053
rect 24213 10013 24225 10047
rect 24259 10013 24271 10047
rect 24213 10007 24271 10013
rect 25961 10047 26019 10053
rect 25961 10013 25973 10047
rect 26007 10044 26019 10047
rect 26234 10044 26240 10056
rect 26007 10016 26240 10044
rect 26007 10013 26019 10016
rect 25961 10007 26019 10013
rect 26234 10004 26240 10016
rect 26292 10004 26298 10056
rect 27264 10053 27292 10152
rect 27614 10072 27620 10124
rect 27672 10072 27678 10124
rect 27893 10115 27951 10121
rect 27893 10081 27905 10115
rect 27939 10112 27951 10115
rect 27982 10112 27988 10124
rect 27939 10084 27988 10112
rect 27939 10081 27951 10084
rect 27893 10075 27951 10081
rect 27982 10072 27988 10084
rect 28040 10072 28046 10124
rect 27249 10047 27307 10053
rect 27249 10013 27261 10047
rect 27295 10044 27307 10047
rect 27295 10016 27660 10044
rect 27295 10013 27307 10016
rect 27249 10007 27307 10013
rect 19245 9979 19303 9985
rect 19245 9945 19257 9979
rect 19291 9976 19303 9979
rect 19720 9976 19748 10004
rect 23201 9979 23259 9985
rect 23201 9976 23213 9979
rect 19291 9948 19748 9976
rect 22112 9948 23213 9976
rect 19291 9945 19303 9948
rect 19245 9939 19303 9945
rect 22112 9917 22140 9948
rect 23201 9945 23213 9948
rect 23247 9945 23259 9979
rect 26252 9976 26280 10004
rect 27632 9988 27660 10016
rect 28994 10004 29000 10056
rect 29052 10004 29058 10056
rect 27341 9979 27399 9985
rect 27341 9976 27353 9979
rect 26252 9948 27353 9976
rect 23201 9939 23259 9945
rect 27341 9945 27353 9948
rect 27387 9945 27399 9979
rect 27341 9939 27399 9945
rect 27525 9979 27583 9985
rect 27525 9945 27537 9979
rect 27571 9945 27583 9979
rect 27525 9939 27583 9945
rect 18064 9880 18828 9908
rect 22097 9911 22155 9917
rect 22097 9877 22109 9911
rect 22143 9877 22155 9911
rect 27540 9908 27568 9939
rect 27614 9936 27620 9988
rect 27672 9936 27678 9988
rect 27798 9908 27804 9920
rect 27540 9880 27804 9908
rect 22097 9871 22155 9877
rect 27798 9868 27804 9880
rect 27856 9908 27862 9920
rect 29365 9911 29423 9917
rect 29365 9908 29377 9911
rect 27856 9880 29377 9908
rect 27856 9868 27862 9880
rect 29365 9877 29377 9880
rect 29411 9877 29423 9911
rect 29365 9871 29423 9877
rect 1104 9818 29716 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 29716 9818
rect 1104 9744 29716 9766
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4856 9676 4905 9704
rect 4856 9664 4862 9676
rect 4893 9673 4905 9676
rect 4939 9673 4951 9707
rect 4893 9667 4951 9673
rect 8849 9707 8907 9713
rect 8849 9673 8861 9707
rect 8895 9704 8907 9707
rect 9030 9704 9036 9716
rect 8895 9676 9036 9704
rect 8895 9673 8907 9676
rect 8849 9667 8907 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 10100 9676 10149 9704
rect 10100 9664 10106 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11422 9704 11428 9716
rect 11020 9676 11428 9704
rect 11020 9664 11026 9676
rect 11422 9664 11428 9676
rect 11480 9704 11486 9716
rect 11480 9676 12020 9704
rect 11480 9664 11486 9676
rect 2130 9596 2136 9648
rect 2188 9596 2194 9648
rect 4522 9596 4528 9648
rect 4580 9636 4586 9648
rect 4985 9639 5043 9645
rect 4985 9636 4997 9639
rect 4580 9608 4997 9636
rect 4580 9596 4586 9608
rect 4985 9605 4997 9608
rect 5031 9636 5043 9639
rect 5994 9636 6000 9648
rect 5031 9608 6000 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5994 9596 6000 9608
rect 6052 9596 6058 9648
rect 7190 9596 7196 9648
rect 7248 9636 7254 9648
rect 7248 9608 7512 9636
rect 7248 9596 7254 9608
rect 3881 9571 3939 9577
rect 3881 9537 3893 9571
rect 3927 9568 3939 9571
rect 4154 9568 4160 9580
rect 3927 9540 4160 9568
rect 3927 9537 3939 9540
rect 3881 9531 3939 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6914 9568 6920 9580
rect 6788 9540 6920 9568
rect 6788 9528 6794 9540
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9566 7159 9571
rect 7208 9566 7236 9596
rect 7484 9577 7512 9608
rect 7147 9538 7236 9566
rect 7377 9571 7435 9577
rect 7147 9537 7159 9538
rect 7101 9531 7159 9537
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9537 7527 9571
rect 7469 9531 7527 9537
rect 8765 9571 8823 9577
rect 8765 9537 8777 9571
rect 8811 9568 8823 9571
rect 9048 9568 9076 9664
rect 9398 9645 9404 9648
rect 9375 9639 9404 9645
rect 9375 9605 9387 9639
rect 9375 9599 9404 9605
rect 9398 9596 9404 9599
rect 9456 9596 9462 9648
rect 11606 9636 11612 9648
rect 9784 9608 11612 9636
rect 9214 9568 9220 9580
rect 9272 9577 9278 9580
rect 9784 9577 9812 9608
rect 11606 9596 11612 9608
rect 11664 9596 11670 9648
rect 11992 9645 12020 9676
rect 13722 9664 13728 9716
rect 13780 9664 13786 9716
rect 17494 9664 17500 9716
rect 17552 9704 17558 9716
rect 18414 9704 18420 9716
rect 17552 9676 18420 9704
rect 17552 9664 17558 9676
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21361 9707 21419 9713
rect 20956 9676 21128 9704
rect 20956 9664 20962 9676
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11955 9608 11989 9636
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13320 9608 13768 9636
rect 13320 9596 13326 9608
rect 13740 9580 13768 9608
rect 14918 9596 14924 9648
rect 14976 9596 14982 9648
rect 21100 9636 21128 9676
rect 21361 9673 21373 9707
rect 21407 9704 21419 9707
rect 21634 9704 21640 9716
rect 21407 9676 21640 9704
rect 21407 9673 21419 9676
rect 21361 9667 21419 9673
rect 21634 9664 21640 9676
rect 21692 9664 21698 9716
rect 21913 9639 21971 9645
rect 21913 9636 21925 9639
rect 21100 9608 21925 9636
rect 9272 9571 9308 9577
rect 8811 9540 8892 9568
rect 9048 9540 9220 9568
rect 8811 9537 8823 9540
rect 8765 9531 8823 9537
rect 1302 9460 1308 9512
rect 1360 9500 1366 9512
rect 1397 9503 1455 9509
rect 1397 9500 1409 9503
rect 1360 9472 1409 9500
rect 1360 9460 1366 9472
rect 1397 9469 1409 9472
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2314 9500 2320 9512
rect 1719 9472 2320 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3421 9503 3479 9509
rect 3421 9500 3433 9503
rect 2740 9472 3433 9500
rect 2740 9460 2746 9472
rect 3421 9469 3433 9472
rect 3467 9469 3479 9503
rect 3421 9463 3479 9469
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 4764 9472 5181 9500
rect 4764 9460 4770 9472
rect 5169 9469 5181 9472
rect 5215 9500 5227 9503
rect 5215 9472 6684 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 6656 9376 6684 9472
rect 6822 9392 6828 9444
rect 6880 9432 6886 9444
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6880 9404 7205 9432
rect 6880 9392 6886 9404
rect 7193 9401 7205 9404
rect 7239 9401 7251 9435
rect 7193 9395 7251 9401
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 2740 9336 3525 9364
rect 2740 9324 2746 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 4614 9364 4620 9376
rect 4571 9336 4620 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 6638 9324 6644 9376
rect 6696 9324 6702 9376
rect 6914 9324 6920 9376
rect 6972 9324 6978 9376
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7392 9364 7420 9531
rect 8864 9512 8892 9540
rect 9214 9528 9220 9540
rect 9296 9537 9308 9571
rect 9272 9531 9308 9537
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 9953 9571 10011 9577
rect 9953 9537 9965 9571
rect 9999 9568 10011 9571
rect 9999 9540 11652 9568
rect 9999 9537 10011 9540
rect 9953 9531 10011 9537
rect 9272 9528 9278 9531
rect 8846 9460 8852 9512
rect 8904 9500 8910 9512
rect 9490 9500 9496 9512
rect 8904 9472 9496 9500
rect 8904 9460 8910 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9582 9460 9588 9512
rect 9640 9460 9646 9512
rect 9674 9460 9680 9512
rect 9732 9492 9738 9512
rect 9876 9492 9904 9531
rect 9732 9464 9904 9492
rect 9732 9460 9738 9464
rect 10134 9460 10140 9512
rect 10192 9460 10198 9512
rect 11624 9509 11652 9540
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 11848 9540 12541 9568
rect 11848 9528 11854 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 13538 9568 13544 9580
rect 12667 9540 13544 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 13633 9571 13691 9577
rect 13633 9537 13645 9571
rect 13679 9537 13691 9571
rect 13633 9531 13691 9537
rect 11609 9503 11667 9509
rect 11609 9469 11621 9503
rect 11655 9500 11667 9503
rect 11882 9500 11888 9512
rect 11655 9472 11888 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 13078 9460 13084 9512
rect 13136 9500 13142 9512
rect 13648 9500 13676 9531
rect 13722 9528 13728 9580
rect 13780 9568 13786 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 13780 9540 13829 9568
rect 13780 9528 13786 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 16666 9568 16672 9580
rect 15059 9540 16672 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17034 9528 17040 9580
rect 17092 9528 17098 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9537 17371 9571
rect 17313 9531 17371 9537
rect 13136 9472 13676 9500
rect 13136 9460 13142 9472
rect 16942 9460 16948 9512
rect 17000 9460 17006 9512
rect 17328 9500 17356 9531
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20312 9540 20913 9568
rect 20312 9528 20318 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9568 21143 9571
rect 21174 9568 21180 9580
rect 21131 9540 21180 9568
rect 21131 9537 21143 9540
rect 21085 9531 21143 9537
rect 19242 9500 19248 9512
rect 17328 9472 19248 9500
rect 19242 9460 19248 9472
rect 19300 9460 19306 9512
rect 9600 9432 9628 9460
rect 9600 9404 9720 9432
rect 7064 9336 7420 9364
rect 9125 9367 9183 9373
rect 7064 9324 7070 9336
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 9582 9364 9588 9376
rect 9171 9336 9588 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9692 9364 9720 9404
rect 10226 9392 10232 9444
rect 10284 9432 10290 9444
rect 12986 9432 12992 9444
rect 10284 9404 12992 9432
rect 10284 9392 10290 9404
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 20916 9432 20944 9531
rect 21174 9528 21180 9540
rect 21232 9528 21238 9580
rect 21468 9577 21496 9608
rect 21913 9605 21925 9608
rect 21959 9605 21971 9639
rect 21913 9599 21971 9605
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22922 9636 22928 9648
rect 22152 9608 22928 9636
rect 22152 9596 22158 9608
rect 22922 9596 22928 9608
rect 22980 9636 22986 9648
rect 23661 9639 23719 9645
rect 23661 9636 23673 9639
rect 22980 9608 23673 9636
rect 22980 9596 22986 9608
rect 23661 9605 23673 9608
rect 23707 9605 23719 9639
rect 23661 9599 23719 9605
rect 23750 9596 23756 9648
rect 23808 9636 23814 9648
rect 24210 9636 24216 9648
rect 23808 9608 24216 9636
rect 23808 9596 23814 9608
rect 24210 9596 24216 9608
rect 24268 9596 24274 9648
rect 26326 9596 26332 9648
rect 26384 9636 26390 9648
rect 27249 9639 27307 9645
rect 27249 9636 27261 9639
rect 26384 9608 27261 9636
rect 26384 9596 26390 9608
rect 27249 9605 27261 9608
rect 27295 9605 27307 9639
rect 27249 9599 27307 9605
rect 27338 9596 27344 9648
rect 27396 9636 27402 9648
rect 27396 9608 27738 9636
rect 27396 9596 27402 9608
rect 28994 9596 29000 9648
rect 29052 9596 29058 9648
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9537 21327 9571
rect 21269 9531 21327 9537
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 20993 9503 21051 9509
rect 20993 9469 21005 9503
rect 21039 9500 21051 9503
rect 21284 9500 21312 9531
rect 21542 9528 21548 9580
rect 21600 9568 21606 9580
rect 21821 9571 21879 9577
rect 21821 9568 21833 9571
rect 21600 9540 21833 9568
rect 21600 9528 21606 9540
rect 21821 9537 21833 9540
rect 21867 9537 21879 9571
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21821 9531 21879 9537
rect 21928 9540 22017 9568
rect 21928 9512 21956 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9537 23535 9571
rect 23477 9531 23535 9537
rect 21039 9472 21312 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 23492 9500 23520 9531
rect 23566 9528 23572 9580
rect 23624 9528 23630 9580
rect 23845 9571 23903 9577
rect 23845 9537 23857 9571
rect 23891 9568 23903 9571
rect 24118 9568 24124 9580
rect 23891 9540 24124 9568
rect 23891 9537 23903 9540
rect 23845 9531 23903 9537
rect 24118 9528 24124 9540
rect 24176 9528 24182 9580
rect 28902 9528 28908 9580
rect 28960 9568 28966 9580
rect 29089 9571 29147 9577
rect 29089 9568 29101 9571
rect 28960 9540 29101 9568
rect 28960 9528 28966 9540
rect 29089 9537 29101 9540
rect 29135 9537 29147 9571
rect 29089 9531 29147 9537
rect 29181 9571 29239 9577
rect 29181 9537 29193 9571
rect 29227 9537 29239 9571
rect 29181 9531 29239 9537
rect 23658 9500 23664 9512
rect 23492 9472 23664 9500
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 25038 9460 25044 9512
rect 25096 9500 25102 9512
rect 26973 9503 27031 9509
rect 26973 9500 26985 9503
rect 25096 9472 26985 9500
rect 25096 9460 25102 9472
rect 26973 9469 26985 9472
rect 27019 9469 27031 9503
rect 26973 9463 27031 9469
rect 27706 9460 27712 9512
rect 27764 9500 27770 9512
rect 28721 9503 28779 9509
rect 28721 9500 28733 9503
rect 27764 9472 28733 9500
rect 27764 9460 27770 9472
rect 28721 9469 28733 9472
rect 28767 9469 28779 9503
rect 28721 9463 28779 9469
rect 21082 9432 21088 9444
rect 20916 9404 21088 9432
rect 21082 9392 21088 9404
rect 21140 9392 21146 9444
rect 26878 9432 26884 9444
rect 22066 9404 26884 9432
rect 11882 9364 11888 9376
rect 9692 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12158 9324 12164 9376
rect 12216 9324 12222 9376
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 15620 9336 16773 9364
rect 15620 9324 15626 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 17497 9367 17555 9373
rect 17497 9333 17509 9367
rect 17543 9364 17555 9367
rect 17586 9364 17592 9376
rect 17543 9336 17592 9364
rect 17543 9333 17555 9336
rect 17497 9327 17555 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 22066 9364 22094 9404
rect 26878 9392 26884 9404
rect 26936 9392 26942 9444
rect 19024 9336 22094 9364
rect 23293 9367 23351 9373
rect 19024 9324 19030 9336
rect 23293 9333 23305 9367
rect 23339 9364 23351 9367
rect 23382 9364 23388 9376
rect 23339 9336 23388 9364
rect 23339 9333 23351 9336
rect 23293 9327 23351 9333
rect 23382 9324 23388 9336
rect 23440 9324 23446 9376
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 29196 9364 29224 9531
rect 29362 9392 29368 9444
rect 29420 9392 29426 9444
rect 24912 9336 29224 9364
rect 24912 9324 24918 9336
rect 1104 9274 29716 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 29716 9274
rect 1104 9200 29716 9222
rect 2130 9120 2136 9172
rect 2188 9120 2194 9172
rect 2314 9120 2320 9172
rect 2372 9120 2378 9172
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 6730 9160 6736 9172
rect 6687 9132 6736 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7558 9160 7564 9172
rect 6840 9132 7564 9160
rect 6840 9092 6868 9132
rect 7558 9120 7564 9132
rect 7616 9160 7622 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 7616 9132 8677 9160
rect 7616 9120 7622 9132
rect 8665 9129 8677 9132
rect 8711 9160 8723 9163
rect 9674 9160 9680 9172
rect 8711 9132 9680 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 9674 9120 9680 9132
rect 9732 9160 9738 9172
rect 10226 9160 10232 9172
rect 9732 9132 10232 9160
rect 9732 9120 9738 9132
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 10643 9132 13124 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 6288 9064 6868 9092
rect 9401 9095 9459 9101
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 2777 9027 2835 9033
rect 2777 9024 2789 9027
rect 2648 8996 2789 9024
rect 2648 8984 2654 8996
rect 2777 8993 2789 8996
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3142 9024 3148 9036
rect 3007 8996 3148 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4614 9024 4620 9036
rect 4295 8996 4620 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2314 8956 2320 8968
rect 2087 8928 2320 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2314 8916 2320 8928
rect 2372 8956 2378 8968
rect 2498 8956 2504 8968
rect 2372 8928 2504 8956
rect 2372 8916 2378 8928
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2682 8916 2688 8968
rect 2740 8916 2746 8968
rect 6288 8965 6316 9064
rect 9401 9061 9413 9095
rect 9447 9092 9459 9095
rect 9447 9064 11284 9092
rect 9447 9061 9459 9064
rect 9401 9055 9459 9061
rect 6362 8984 6368 9036
rect 6420 8984 6426 9036
rect 8846 9024 8852 9036
rect 6748 8996 8852 9024
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 3988 8820 4016 8919
rect 5258 8848 5264 8900
rect 5316 8848 5322 8900
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6748 8888 6776 8996
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9088 8996 9168 9024
rect 9088 8984 9094 8996
rect 9140 8965 9168 8996
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9640 8996 9873 9024
rect 9640 8984 9646 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10091 8996 11192 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6052 8860 6776 8888
rect 6840 8928 6929 8956
rect 6840 8888 6868 8928
rect 6917 8925 6929 8928
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 7098 8888 7104 8900
rect 6840 8860 7104 8888
rect 6052 8848 6058 8860
rect 6454 8820 6460 8832
rect 3988 8792 6460 8820
rect 6454 8780 6460 8792
rect 6512 8820 6518 8832
rect 6840 8820 6868 8860
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7190 8848 7196 8900
rect 7248 8848 7254 8900
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 8418 8860 9045 8888
rect 9033 8857 9045 8860
rect 9079 8857 9091 8891
rect 9876 8888 9904 8987
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10376 8928 10425 8956
rect 10376 8916 10382 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10502 8916 10508 8968
rect 10560 8916 10566 8968
rect 11164 8965 11192 8996
rect 10781 8959 10839 8965
rect 10781 8956 10793 8959
rect 10612 8928 10793 8956
rect 10612 8888 10640 8928
rect 10781 8925 10793 8928
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8925 11115 8959
rect 11057 8919 11115 8925
rect 11150 8959 11208 8965
rect 11150 8925 11162 8959
rect 11196 8925 11208 8959
rect 11150 8919 11208 8925
rect 9876 8860 10640 8888
rect 10689 8891 10747 8897
rect 9033 8851 9091 8857
rect 10689 8857 10701 8891
rect 10735 8888 10747 8891
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10735 8860 10885 8888
rect 10735 8857 10747 8860
rect 10689 8851 10747 8857
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 11072 8888 11100 8919
rect 11256 8900 11284 9064
rect 12158 8984 12164 9036
rect 12216 9024 12222 9036
rect 12216 8996 12664 9024
rect 12216 8984 12222 8996
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11563 8959 11621 8965
rect 11563 8925 11575 8959
rect 11609 8956 11621 8959
rect 11790 8956 11796 8968
rect 11609 8928 11796 8956
rect 11609 8925 11621 8928
rect 11563 8919 11621 8925
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 12636 8965 12664 8996
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8925 12679 8959
rect 12621 8919 12679 8925
rect 11238 8888 11244 8900
rect 11072 8860 11244 8888
rect 10873 8851 10931 8857
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8857 11391 8891
rect 12360 8888 12388 8919
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 12894 8916 12900 8968
rect 12952 8916 12958 8968
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 13096 8956 13124 9132
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 13228 9132 13369 9160
rect 13228 9120 13234 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 16942 9120 16948 9172
rect 17000 9120 17006 9172
rect 22002 9160 22008 9172
rect 17236 9132 22008 9160
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13311 8996 13645 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 13725 9027 13783 9033
rect 13725 8993 13737 9027
rect 13771 9024 13783 9027
rect 15654 9024 15660 9036
rect 13771 8996 15660 9024
rect 13771 8993 13783 8996
rect 13725 8987 13783 8993
rect 15654 8984 15660 8996
rect 15712 8984 15718 9036
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 9024 15899 9027
rect 16390 9024 16396 9036
rect 15887 8996 16396 9024
rect 15887 8993 15899 8996
rect 15841 8987 15899 8993
rect 16390 8984 16396 8996
rect 16448 8984 16454 9036
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 13096 8928 13553 8956
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13817 8959 13875 8965
rect 13817 8925 13829 8959
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 11333 8851 11391 8857
rect 11716 8860 12388 8888
rect 12529 8891 12587 8897
rect 6512 8792 6868 8820
rect 6512 8780 6518 8792
rect 10226 8780 10232 8832
rect 10284 8780 10290 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 11348 8820 11376 8851
rect 11716 8829 11744 8860
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 13832 8888 13860 8919
rect 15562 8916 15568 8968
rect 15620 8916 15626 8968
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 17092 8928 17141 8956
rect 17092 8916 17098 8928
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17236 8888 17264 9132
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23017 9163 23075 9169
rect 23017 9160 23029 9163
rect 22152 9132 23029 9160
rect 22152 9120 22158 9132
rect 23017 9129 23029 9132
rect 23063 9129 23075 9163
rect 23017 9123 23075 9129
rect 27338 9120 27344 9172
rect 27396 9120 27402 9172
rect 19242 9052 19248 9104
rect 19300 9052 19306 9104
rect 22186 9052 22192 9104
rect 22244 9092 22250 9104
rect 22373 9095 22431 9101
rect 22373 9092 22385 9095
rect 22244 9064 22385 9092
rect 22244 9052 22250 9064
rect 22373 9061 22385 9064
rect 22419 9061 22431 9095
rect 22373 9055 22431 9061
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17420 8996 17785 9024
rect 17420 8968 17448 8996
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 20993 9027 21051 9033
rect 20993 9024 21005 9027
rect 20772 8996 21005 9024
rect 20772 8984 20778 8996
rect 20993 8993 21005 8996
rect 21039 8993 21051 9027
rect 23106 9024 23112 9036
rect 20993 8987 21051 8993
rect 22112 8996 23112 9024
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17586 8916 17592 8968
rect 17644 8916 17650 8968
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 21082 8916 21088 8968
rect 21140 8956 21146 8968
rect 22112 8965 22140 8996
rect 23106 8984 23112 8996
rect 23164 8984 23170 9036
rect 23308 8996 23888 9024
rect 22097 8959 22155 8965
rect 22097 8956 22109 8959
rect 21140 8928 22109 8956
rect 21140 8916 21146 8928
rect 22097 8925 22109 8928
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22370 8916 22376 8968
rect 22428 8956 22434 8968
rect 22649 8959 22707 8965
rect 22649 8956 22661 8959
rect 22428 8928 22661 8956
rect 22428 8916 22434 8928
rect 22649 8925 22661 8928
rect 22695 8925 22707 8959
rect 22649 8919 22707 8925
rect 23196 8959 23254 8965
rect 23196 8925 23208 8959
rect 23242 8956 23254 8959
rect 23308 8956 23336 8996
rect 23242 8928 23336 8956
rect 23242 8925 23254 8928
rect 23196 8919 23254 8925
rect 23382 8916 23388 8968
rect 23440 8916 23446 8968
rect 23474 8916 23480 8968
rect 23532 8965 23538 8968
rect 23532 8959 23571 8965
rect 23559 8925 23571 8959
rect 23532 8919 23571 8925
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8925 23719 8959
rect 23661 8919 23719 8925
rect 23532 8916 23538 8919
rect 12575 8860 13860 8888
rect 14660 8860 17264 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 10560 8792 11376 8820
rect 11701 8823 11759 8829
rect 10560 8780 10566 8792
rect 11701 8789 11713 8823
rect 11747 8789 11759 8823
rect 11701 8783 11759 8789
rect 11882 8780 11888 8832
rect 11940 8820 11946 8832
rect 14660 8820 14688 8860
rect 20070 8848 20076 8900
rect 20128 8848 20134 8900
rect 20717 8891 20775 8897
rect 20717 8857 20729 8891
rect 20763 8857 20775 8891
rect 20717 8851 20775 8857
rect 22741 8891 22799 8897
rect 22741 8857 22753 8891
rect 22787 8888 22799 8891
rect 23290 8888 23296 8900
rect 22787 8860 23296 8888
rect 22787 8857 22799 8860
rect 22741 8851 22799 8857
rect 11940 8792 14688 8820
rect 11940 8780 11946 8792
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 14792 8792 15209 8820
rect 14792 8780 14798 8792
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 15197 8783 15255 8789
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 16206 8820 16212 8832
rect 15703 8792 16212 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 16206 8780 16212 8792
rect 16264 8780 16270 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17678 8820 17684 8832
rect 16724 8792 17684 8820
rect 16724 8780 16730 8792
rect 17678 8780 17684 8792
rect 17736 8780 17742 8832
rect 18230 8780 18236 8832
rect 18288 8780 18294 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 20732 8820 20760 8851
rect 23290 8848 23296 8860
rect 23348 8848 23354 8900
rect 23676 8888 23704 8919
rect 23860 8900 23888 8996
rect 24486 8916 24492 8968
rect 24544 8916 24550 8968
rect 26418 8916 26424 8968
rect 26476 8956 26482 8968
rect 27249 8959 27307 8965
rect 27249 8956 27261 8959
rect 26476 8928 27261 8956
rect 26476 8916 26482 8928
rect 27249 8925 27261 8928
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 23492 8860 23704 8888
rect 19760 8792 20760 8820
rect 19760 8780 19766 8792
rect 20898 8780 20904 8832
rect 20956 8820 20962 8832
rect 21177 8823 21235 8829
rect 21177 8820 21189 8823
rect 20956 8792 21189 8820
rect 20956 8780 20962 8792
rect 21177 8789 21189 8792
rect 21223 8789 21235 8823
rect 21177 8783 21235 8789
rect 22557 8823 22615 8829
rect 22557 8789 22569 8823
rect 22603 8820 22615 8823
rect 23492 8820 23520 8860
rect 23842 8848 23848 8900
rect 23900 8888 23906 8900
rect 28626 8888 28632 8900
rect 23900 8860 28632 8888
rect 23900 8848 23906 8860
rect 28626 8848 28632 8860
rect 28684 8848 28690 8900
rect 22603 8792 23520 8820
rect 22603 8789 22615 8792
rect 22557 8783 22615 8789
rect 23566 8780 23572 8832
rect 23624 8820 23630 8832
rect 24581 8823 24639 8829
rect 24581 8820 24593 8823
rect 23624 8792 24593 8820
rect 23624 8780 23630 8792
rect 24581 8789 24593 8792
rect 24627 8820 24639 8823
rect 24670 8820 24676 8832
rect 24627 8792 24676 8820
rect 24627 8789 24639 8792
rect 24581 8783 24639 8789
rect 24670 8780 24676 8792
rect 24728 8780 24734 8832
rect 1104 8730 29716 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 29716 8730
rect 1104 8656 29716 8678
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5258 8616 5264 8628
rect 5123 8588 5264 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 7190 8616 7196 8628
rect 6963 8588 7196 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 9122 8616 9128 8628
rect 7300 8588 9128 8616
rect 7300 8548 7328 8588
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 11606 8576 11612 8628
rect 11664 8576 11670 8628
rect 12627 8619 12685 8625
rect 12627 8585 12639 8619
rect 12673 8616 12685 8619
rect 12802 8616 12808 8628
rect 12673 8588 12808 8616
rect 12673 8585 12685 8588
rect 12627 8579 12685 8585
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13872 8588 13921 8616
rect 13872 8576 13878 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 16206 8576 16212 8628
rect 16264 8616 16270 8628
rect 16264 8588 16528 8616
rect 16264 8576 16270 8588
rect 1688 8520 7328 8548
rect 1688 8489 1716 8520
rect 7558 8508 7564 8560
rect 7616 8508 7622 8560
rect 11238 8508 11244 8560
rect 11296 8548 11302 8560
rect 12529 8551 12587 8557
rect 12529 8548 12541 8551
rect 11296 8520 12541 8548
rect 11296 8508 11302 8520
rect 12529 8517 12541 8520
rect 12575 8517 12587 8551
rect 12529 8511 12587 8517
rect 14734 8508 14740 8560
rect 14792 8508 14798 8560
rect 15470 8508 15476 8560
rect 15528 8508 15534 8560
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 16393 8551 16451 8557
rect 16393 8548 16405 8551
rect 16172 8520 16405 8548
rect 16172 8508 16178 8520
rect 16393 8517 16405 8520
rect 16439 8517 16451 8551
rect 16393 8511 16451 8517
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 2372 8452 4997 8480
rect 2372 8440 2378 8452
rect 4985 8449 4997 8452
rect 5031 8480 5043 8483
rect 5626 8480 5632 8492
rect 5031 8452 5632 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 6972 8452 7205 8480
rect 6972 8440 6978 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 12342 8480 12348 8492
rect 11747 8452 12348 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 12434 8440 12440 8492
rect 12492 8480 12498 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12492 8452 12725 8480
rect 12492 8440 12498 8452
rect 12713 8449 12725 8452
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 12986 8480 12992 8492
rect 12851 8452 12992 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13814 8440 13820 8492
rect 13872 8440 13878 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6880 8384 7113 8412
rect 6880 8372 6886 8384
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7466 8372 7472 8424
rect 7524 8372 7530 8424
rect 9398 8372 9404 8424
rect 9456 8412 9462 8424
rect 12526 8412 12532 8424
rect 9456 8384 12532 8412
rect 9456 8372 9462 8384
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 13446 8372 13452 8424
rect 13504 8412 13510 8424
rect 13722 8412 13728 8424
rect 13504 8384 13728 8412
rect 13504 8372 13510 8384
rect 13722 8372 13728 8384
rect 13780 8412 13786 8424
rect 14016 8412 14044 8443
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 16500 8489 16528 8588
rect 17034 8576 17040 8628
rect 17092 8576 17098 8628
rect 17405 8619 17463 8625
rect 17405 8585 17417 8619
rect 17451 8616 17463 8619
rect 17862 8616 17868 8628
rect 17451 8588 17868 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 19245 8619 19303 8625
rect 19245 8616 19257 8619
rect 18288 8588 19257 8616
rect 18288 8576 18294 8588
rect 19245 8585 19257 8588
rect 19291 8585 19303 8619
rect 19245 8579 19303 8585
rect 19613 8619 19671 8625
rect 19613 8585 19625 8619
rect 19659 8616 19671 8619
rect 19702 8616 19708 8628
rect 19659 8588 19708 8616
rect 19659 8585 19671 8588
rect 19613 8579 19671 8585
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20070 8576 20076 8628
rect 20128 8576 20134 8628
rect 23385 8619 23443 8625
rect 23385 8585 23397 8619
rect 23431 8616 23443 8619
rect 23474 8616 23480 8628
rect 23431 8588 23480 8616
rect 23431 8585 23443 8588
rect 23385 8579 23443 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 23658 8576 23664 8628
rect 23716 8576 23722 8628
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24946 8616 24952 8628
rect 24176 8588 24952 8616
rect 24176 8576 24182 8588
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 26878 8576 26884 8628
rect 26936 8616 26942 8628
rect 29181 8619 29239 8625
rect 29181 8616 29193 8619
rect 26936 8588 29193 8616
rect 26936 8576 26942 8588
rect 29181 8585 29193 8588
rect 29227 8585 29239 8619
rect 29181 8579 29239 8585
rect 17052 8548 17080 8576
rect 17052 8520 17356 8548
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14332 8452 14473 8480
rect 14332 8440 14338 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8480 17003 8483
rect 17034 8480 17040 8492
rect 16991 8452 17040 8480
rect 16991 8449 17003 8452
rect 16945 8443 17003 8449
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17218 8480 17224 8492
rect 17175 8452 17224 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 17328 8489 17356 8520
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 22186 8548 22192 8560
rect 17736 8520 20208 8548
rect 17736 8508 17742 8520
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8449 17371 8483
rect 17313 8443 17371 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17586 8480 17592 8492
rect 17543 8452 17592 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 19153 8483 19211 8489
rect 19153 8449 19165 8483
rect 19199 8480 19211 8483
rect 19242 8480 19248 8492
rect 19199 8452 19248 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 20180 8489 20208 8520
rect 20272 8520 22192 8548
rect 20272 8492 20300 8520
rect 22186 8508 22192 8520
rect 22244 8508 22250 8560
rect 23676 8548 23704 8576
rect 23584 8520 23704 8548
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 20254 8440 20260 8492
rect 20312 8440 20318 8492
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 20622 8480 20628 8492
rect 20404 8452 20628 8480
rect 20404 8440 20410 8452
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 23474 8480 23480 8492
rect 22066 8452 23480 8480
rect 13780 8384 14044 8412
rect 14568 8384 15792 8412
rect 13780 8372 13786 8384
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 14568 8344 14596 8384
rect 2464 8316 14596 8344
rect 15764 8344 15792 8384
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 18969 8415 19027 8421
rect 18969 8412 18981 8415
rect 16448 8384 18981 8412
rect 16448 8372 16454 8384
rect 18969 8381 18981 8384
rect 19015 8381 19027 8415
rect 18969 8375 19027 8381
rect 22066 8344 22094 8452
rect 23474 8440 23480 8452
rect 23532 8480 23538 8492
rect 23584 8489 23612 8520
rect 23569 8483 23627 8489
rect 23569 8480 23581 8483
rect 23532 8452 23581 8480
rect 23532 8440 23538 8452
rect 23569 8449 23581 8452
rect 23615 8449 23627 8483
rect 23569 8443 23627 8449
rect 23658 8440 23664 8492
rect 23716 8440 23722 8492
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 23290 8372 23296 8424
rect 23348 8412 23354 8424
rect 23952 8412 23980 8443
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8480 25743 8483
rect 28166 8480 28172 8492
rect 25731 8452 28172 8480
rect 25731 8449 25743 8452
rect 25685 8443 25743 8449
rect 28166 8440 28172 8452
rect 28224 8440 28230 8492
rect 29270 8440 29276 8492
rect 29328 8440 29334 8492
rect 23348 8384 23980 8412
rect 23348 8372 23354 8384
rect 15764 8316 22094 8344
rect 2464 8304 2470 8316
rect 23842 8304 23848 8356
rect 23900 8304 23906 8356
rect 24118 8304 24124 8356
rect 24176 8344 24182 8356
rect 25593 8347 25651 8353
rect 25593 8344 25605 8347
rect 24176 8316 25605 8344
rect 24176 8304 24182 8316
rect 25593 8313 25605 8316
rect 25639 8313 25651 8347
rect 25593 8307 25651 8313
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 8018 8276 8024 8288
rect 1820 8248 8024 8276
rect 1820 8236 1826 8248
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 10962 8276 10968 8288
rect 9916 8248 10968 8276
rect 9916 8236 9922 8248
rect 10962 8236 10968 8248
rect 11020 8236 11026 8288
rect 11606 8236 11612 8288
rect 11664 8276 11670 8288
rect 12434 8276 12440 8288
rect 11664 8248 12440 8276
rect 11664 8236 11670 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 20441 8279 20499 8285
rect 20441 8245 20453 8279
rect 20487 8276 20499 8279
rect 20530 8276 20536 8288
rect 20487 8248 20536 8276
rect 20487 8245 20499 8248
rect 20441 8239 20499 8245
rect 20530 8236 20536 8248
rect 20588 8236 20594 8288
rect 20898 8236 20904 8288
rect 20956 8276 20962 8288
rect 21910 8276 21916 8288
rect 20956 8248 21916 8276
rect 20956 8236 20962 8248
rect 21910 8236 21916 8248
rect 21968 8276 21974 8288
rect 23382 8276 23388 8288
rect 21968 8248 23388 8276
rect 21968 8236 21974 8248
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 1104 8186 29716 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 29716 8186
rect 1104 8112 29716 8134
rect 6273 8075 6331 8081
rect 2746 8044 6224 8072
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2746 7936 2774 8044
rect 3068 7976 3464 8004
rect 3068 7945 3096 7976
rect 1719 7908 2774 7936
rect 3053 7939 3111 7945
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 3053 7905 3065 7939
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7905 3387 7939
rect 3436 7936 3464 7976
rect 4706 7964 4712 8016
rect 4764 8004 4770 8016
rect 6196 8004 6224 8044
rect 6273 8041 6285 8075
rect 6319 8072 6331 8075
rect 7282 8072 7288 8084
rect 6319 8044 7288 8072
rect 6319 8041 6331 8044
rect 6273 8035 6331 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 10318 8032 10324 8084
rect 10376 8032 10382 8084
rect 11425 8075 11483 8081
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 11698 8072 11704 8084
rect 11471 8044 11704 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12253 8075 12311 8081
rect 12253 8041 12265 8075
rect 12299 8072 12311 8075
rect 12618 8072 12624 8084
rect 12299 8044 12624 8072
rect 12299 8041 12311 8044
rect 12253 8035 12311 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13814 8032 13820 8084
rect 13872 8032 13878 8084
rect 15470 8032 15476 8084
rect 15528 8072 15534 8084
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 15528 8044 15577 8072
rect 15528 8032 15534 8044
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 15565 8035 15623 8041
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 22278 8072 22284 8084
rect 21324 8044 22284 8072
rect 21324 8032 21330 8044
rect 22278 8032 22284 8044
rect 22336 8072 22342 8084
rect 22336 8044 22784 8072
rect 22336 8032 22342 8044
rect 9398 8004 9404 8016
rect 4764 7976 6040 8004
rect 6196 7976 9404 8004
rect 4764 7964 4770 7976
rect 4798 7936 4804 7948
rect 3436 7908 4804 7936
rect 3329 7899 3387 7905
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 2958 7828 2964 7880
rect 3016 7828 3022 7880
rect 3344 7800 3372 7899
rect 4798 7896 4804 7908
rect 4856 7936 4862 7948
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4856 7908 4997 7936
rect 4856 7896 4862 7908
rect 4985 7905 4997 7908
rect 5031 7905 5043 7939
rect 5810 7936 5816 7948
rect 4985 7899 5043 7905
rect 5092 7908 5816 7936
rect 5092 7877 5120 7908
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 5902 7896 5908 7948
rect 5960 7896 5966 7948
rect 6012 7945 6040 7976
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 10962 7964 10968 8016
rect 11020 7964 11026 8016
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 11112 7976 11560 8004
rect 11112 7964 11118 7976
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 5997 7899 6055 7905
rect 6748 7908 9689 7936
rect 5077 7871 5135 7877
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 5718 7868 5724 7880
rect 5675 7840 5724 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 5718 7828 5724 7840
rect 5776 7868 5782 7880
rect 6748 7868 6776 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 11072 7908 11284 7936
rect 5776 7840 6776 7868
rect 5776 7828 5782 7840
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7101 7871 7159 7877
rect 7101 7868 7113 7871
rect 6932 7840 7113 7868
rect 4430 7800 4436 7812
rect 3344 7772 4436 7800
rect 4430 7760 4436 7772
rect 4488 7800 4494 7812
rect 6114 7803 6172 7809
rect 6114 7800 6126 7803
rect 4488 7772 6126 7800
rect 4488 7760 4494 7772
rect 6114 7769 6126 7772
rect 6160 7769 6172 7803
rect 6114 7763 6172 7769
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 6932 7800 6960 7840
rect 7101 7837 7113 7840
rect 7147 7868 7159 7871
rect 7282 7868 7288 7880
rect 7147 7840 7288 7868
rect 7147 7837 7159 7840
rect 7101 7831 7159 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 8076 7840 8125 7868
rect 8076 7828 8082 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 6420 7772 6960 7800
rect 7009 7803 7067 7809
rect 6420 7760 6426 7772
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 7558 7800 7564 7812
rect 7055 7772 7564 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 6380 7732 6408 7760
rect 7116 7744 7144 7772
rect 7558 7760 7564 7772
rect 7616 7760 7622 7812
rect 8128 7800 8156 7831
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9548 7840 9597 7868
rect 9548 7828 9554 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7868 9827 7871
rect 10042 7868 10048 7880
rect 9815 7840 10048 7868
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10318 7828 10324 7880
rect 10376 7868 10382 7880
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10376 7840 10517 7868
rect 10376 7828 10382 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 10643 7840 10824 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 8478 7800 8484 7812
rect 8128 7772 8484 7800
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 10612 7800 10640 7831
rect 10468 7772 10640 7800
rect 10689 7803 10747 7809
rect 10468 7760 10474 7772
rect 10689 7769 10701 7803
rect 10735 7769 10747 7803
rect 10796 7800 10824 7840
rect 10870 7828 10876 7880
rect 10928 7828 10934 7880
rect 11072 7868 11100 7908
rect 10980 7840 11100 7868
rect 10980 7800 11008 7840
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 11256 7877 11284 7908
rect 11532 7877 11560 7976
rect 13556 7976 14504 8004
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 13556 7936 13584 7976
rect 13814 7936 13820 7948
rect 11756 7908 13584 7936
rect 13648 7908 13820 7936
rect 11756 7896 11762 7908
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11790 7828 11796 7880
rect 11848 7868 11854 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11848 7840 11897 7868
rect 11848 7828 11854 7840
rect 11885 7837 11897 7840
rect 11931 7868 11943 7871
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 11931 7840 13001 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7868 13139 7871
rect 13446 7868 13452 7880
rect 13127 7840 13452 7868
rect 13127 7837 13139 7840
rect 13081 7831 13139 7837
rect 13446 7828 13452 7840
rect 13504 7828 13510 7880
rect 13648 7877 13676 7908
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 14476 7880 14504 7976
rect 19812 7976 21495 8004
rect 19812 7936 19840 7976
rect 19720 7908 19840 7936
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13964 7840 14105 7868
rect 13964 7828 13970 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 14277 7871 14335 7877
rect 14277 7868 14289 7871
rect 14240 7840 14289 7868
rect 14240 7828 14246 7840
rect 14277 7837 14289 7840
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 14366 7828 14372 7880
rect 14424 7828 14430 7880
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 15473 7871 15531 7877
rect 15473 7837 15485 7871
rect 15519 7868 15531 7871
rect 16666 7868 16672 7880
rect 15519 7840 16672 7868
rect 15519 7837 15531 7840
rect 15473 7831 15531 7837
rect 16666 7828 16672 7840
rect 16724 7828 16730 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 18046 7868 18052 7880
rect 17267 7840 18052 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 18046 7828 18052 7840
rect 18104 7868 18110 7880
rect 19242 7868 19248 7880
rect 18104 7840 19248 7868
rect 18104 7828 18110 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19720 7877 19748 7908
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20162 7936 20168 7948
rect 19944 7908 20168 7936
rect 19944 7896 19950 7908
rect 20162 7896 20168 7908
rect 20220 7936 20226 7948
rect 20220 7908 20484 7936
rect 20220 7896 20226 7908
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19392 7840 19533 7868
rect 19392 7828 19398 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7837 19763 7871
rect 19705 7831 19763 7837
rect 19797 7871 19855 7877
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 20070 7868 20076 7880
rect 19843 7840 20076 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20456 7877 20484 7908
rect 20622 7896 20628 7948
rect 20680 7936 20686 7948
rect 20680 7908 20944 7936
rect 20680 7896 20686 7908
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 10796 7772 11008 7800
rect 10689 7763 10747 7769
rect 6052 7704 6408 7732
rect 6052 7692 6058 7704
rect 6638 7692 6644 7744
rect 6696 7692 6702 7744
rect 7098 7692 7104 7744
rect 7156 7692 7162 7744
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 8021 7735 8079 7741
rect 8021 7732 8033 7735
rect 7984 7704 8033 7732
rect 7984 7692 7990 7704
rect 8021 7701 8033 7704
rect 8067 7701 8079 7735
rect 8021 7695 8079 7701
rect 8294 7692 8300 7744
rect 8352 7692 8358 7744
rect 10704 7732 10732 7763
rect 12066 7760 12072 7812
rect 12124 7760 12130 7812
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 14829 7803 14887 7809
rect 14829 7800 14841 7803
rect 12216 7772 14841 7800
rect 12216 7760 12222 7772
rect 14829 7769 14841 7772
rect 14875 7769 14887 7803
rect 14829 7763 14887 7769
rect 19978 7760 19984 7812
rect 20036 7800 20042 7812
rect 20364 7800 20392 7831
rect 20530 7828 20536 7880
rect 20588 7828 20594 7880
rect 20916 7877 20944 7908
rect 20990 7896 20996 7948
rect 21048 7896 21054 7948
rect 21467 7936 21495 7976
rect 21818 7964 21824 8016
rect 21876 7964 21882 8016
rect 22005 8007 22063 8013
rect 22005 7973 22017 8007
rect 22051 8004 22063 8007
rect 22646 8004 22652 8016
rect 22051 7976 22652 8004
rect 22051 7973 22063 7976
rect 22005 7967 22063 7973
rect 22646 7964 22652 7976
rect 22704 7964 22710 8016
rect 22756 8004 22784 8044
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 24026 8072 24032 8084
rect 22888 8044 24032 8072
rect 22888 8032 22894 8044
rect 24026 8032 24032 8044
rect 24084 8032 24090 8084
rect 24118 8032 24124 8084
rect 24176 8032 24182 8084
rect 24136 8004 24164 8032
rect 22756 7976 24164 8004
rect 22554 7936 22560 7948
rect 21100 7908 21404 7936
rect 21467 7908 22560 7936
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 20036 7772 20392 7800
rect 20732 7800 20760 7831
rect 21100 7800 21128 7908
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 20732 7772 21128 7800
rect 20036 7760 20042 7772
rect 11054 7732 11060 7744
rect 10704 7704 11060 7732
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 13538 7692 13544 7744
rect 13596 7692 13602 7744
rect 17126 7692 17132 7744
rect 17184 7732 17190 7744
rect 17678 7732 17684 7744
rect 17184 7704 17684 7732
rect 17184 7692 17190 7704
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 19426 7732 19432 7744
rect 19383 7704 19432 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 20162 7692 20168 7744
rect 20220 7692 20226 7744
rect 21192 7732 21220 7831
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 21376 7868 21404 7908
rect 22554 7896 22560 7908
rect 22612 7896 22618 7948
rect 23753 7939 23811 7945
rect 23753 7936 23765 7939
rect 22848 7908 23765 7936
rect 22094 7868 22100 7880
rect 21376 7840 22100 7868
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 22278 7877 22284 7880
rect 22276 7868 22284 7877
rect 22239 7840 22284 7868
rect 22276 7831 22284 7840
rect 22278 7828 22284 7831
rect 22336 7828 22342 7880
rect 22370 7828 22376 7880
rect 22428 7828 22434 7880
rect 22646 7868 22652 7880
rect 22607 7840 22652 7868
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 22738 7828 22744 7880
rect 22796 7828 22802 7880
rect 21450 7760 21456 7812
rect 21508 7760 21514 7812
rect 21542 7760 21548 7812
rect 21600 7760 21606 7812
rect 22388 7800 22416 7828
rect 21652 7772 22416 7800
rect 22465 7803 22523 7809
rect 21652 7732 21680 7772
rect 22465 7769 22477 7803
rect 22511 7769 22523 7803
rect 22465 7763 22523 7769
rect 21192 7704 21680 7732
rect 22094 7692 22100 7744
rect 22152 7692 22158 7744
rect 22278 7692 22284 7744
rect 22336 7732 22342 7744
rect 22480 7732 22508 7763
rect 22554 7760 22560 7812
rect 22612 7800 22618 7812
rect 22848 7800 22876 7908
rect 23753 7905 23765 7908
rect 23799 7905 23811 7939
rect 29546 7936 29552 7948
rect 23753 7899 23811 7905
rect 24596 7908 29552 7936
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23198 7868 23204 7880
rect 23155 7840 23204 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 23382 7828 23388 7880
rect 23440 7828 23446 7880
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7837 23995 7871
rect 23937 7831 23995 7837
rect 22612 7772 22876 7800
rect 23293 7803 23351 7809
rect 22612 7760 22618 7772
rect 23293 7769 23305 7803
rect 23339 7800 23351 7803
rect 23842 7800 23848 7812
rect 23339 7772 23848 7800
rect 23339 7769 23351 7772
rect 23293 7763 23351 7769
rect 23842 7760 23848 7772
rect 23900 7760 23906 7812
rect 22336 7704 22508 7732
rect 23661 7735 23719 7741
rect 22336 7692 22342 7704
rect 23661 7701 23673 7735
rect 23707 7732 23719 7735
rect 23952 7732 23980 7831
rect 24210 7828 24216 7880
rect 24268 7828 24274 7880
rect 24394 7828 24400 7880
rect 24452 7868 24458 7880
rect 24596 7877 24624 7908
rect 29546 7896 29552 7908
rect 29604 7896 29610 7948
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 24452 7840 24593 7868
rect 24452 7828 24458 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 24670 7828 24676 7880
rect 24728 7828 24734 7880
rect 24946 7828 24952 7880
rect 25004 7828 25010 7880
rect 29362 7828 29368 7880
rect 29420 7828 29426 7880
rect 24302 7760 24308 7812
rect 24360 7800 24366 7812
rect 24765 7803 24823 7809
rect 24765 7800 24777 7803
rect 24360 7772 24777 7800
rect 24360 7760 24366 7772
rect 24765 7769 24777 7772
rect 24811 7800 24823 7803
rect 29730 7800 29736 7812
rect 24811 7772 29736 7800
rect 24811 7769 24823 7772
rect 24765 7763 24823 7769
rect 29730 7760 29736 7772
rect 29788 7760 29794 7812
rect 23707 7704 23980 7732
rect 24121 7735 24179 7741
rect 23707 7701 23719 7704
rect 23661 7695 23719 7701
rect 24121 7701 24133 7735
rect 24167 7732 24179 7735
rect 24397 7735 24455 7741
rect 24397 7732 24409 7735
rect 24167 7704 24409 7732
rect 24167 7701 24179 7704
rect 24121 7695 24179 7701
rect 24397 7701 24409 7704
rect 24443 7701 24455 7735
rect 24397 7695 24455 7701
rect 29178 7692 29184 7744
rect 29236 7692 29242 7744
rect 1104 7642 29716 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 29716 7642
rect 1104 7568 29716 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 2915 7500 3341 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6641 7531 6699 7537
rect 6641 7528 6653 7531
rect 6604 7500 6653 7528
rect 6604 7488 6610 7500
rect 6641 7497 6653 7500
rect 6687 7497 6699 7531
rect 6641 7491 6699 7497
rect 8202 7488 8208 7540
rect 8260 7488 8266 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 10410 7528 10416 7540
rect 8352 7500 10416 7528
rect 8352 7488 8358 7500
rect 4065 7463 4123 7469
rect 4065 7460 4077 7463
rect 3804 7432 4077 7460
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 2958 7284 2964 7336
rect 3016 7284 3022 7336
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 1670 7148 1676 7200
rect 1728 7188 1734 7200
rect 2501 7191 2559 7197
rect 2501 7188 2513 7191
rect 1728 7160 2513 7188
rect 1728 7148 1734 7160
rect 2501 7157 2513 7160
rect 2547 7157 2559 7191
rect 2976 7188 3004 7284
rect 3712 7256 3740 7355
rect 3804 7333 3832 7432
rect 4065 7429 4077 7432
rect 4111 7460 4123 7463
rect 5445 7463 5503 7469
rect 5445 7460 5457 7463
rect 4111 7432 5457 7460
rect 4111 7429 4123 7432
rect 4065 7423 4123 7429
rect 5445 7429 5457 7432
rect 5491 7429 5503 7463
rect 6086 7460 6092 7472
rect 5445 7423 5503 7429
rect 5552 7432 6092 7460
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4632 7324 4660 7355
rect 4571 7296 4660 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4430 7256 4436 7268
rect 3712 7228 4436 7256
rect 4430 7216 4436 7228
rect 4488 7216 4494 7268
rect 4816 7256 4844 7355
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 4540 7228 4844 7256
rect 4908 7256 4936 7352
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 5552 7324 5580 7432
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 5982 7401 6010 7432
rect 6086 7420 6092 7432
rect 6144 7460 6150 7472
rect 7193 7463 7251 7469
rect 7193 7460 7205 7463
rect 6144 7432 7205 7460
rect 6144 7420 6150 7432
rect 7193 7429 7205 7432
rect 7239 7429 7251 7463
rect 7193 7423 7251 7429
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 7561 7463 7619 7469
rect 7561 7460 7573 7463
rect 7340 7432 7573 7460
rect 7340 7420 7346 7432
rect 7561 7429 7573 7432
rect 7607 7429 7619 7463
rect 8220 7460 8248 7488
rect 7561 7423 7619 7429
rect 8036 7432 8248 7460
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5776 7364 5825 7392
rect 5776 7352 5782 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5967 7395 6025 7401
rect 5967 7361 5979 7395
rect 6013 7361 6025 7395
rect 5967 7355 6025 7361
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6822 7392 6828 7404
rect 6236 7364 6828 7392
rect 6236 7352 6242 7364
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7926 7352 7932 7404
rect 7984 7352 7990 7404
rect 8036 7401 8064 7432
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 5491 7296 5580 7324
rect 5629 7327 5687 7333
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 6638 7324 6644 7336
rect 5675 7296 6644 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7392 7324 7420 7352
rect 7055 7296 7420 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 5994 7256 6000 7268
rect 4908 7228 6000 7256
rect 4540 7188 4568 7228
rect 2976 7160 4568 7188
rect 2501 7151 2559 7157
rect 4614 7148 4620 7200
rect 4672 7148 4678 7200
rect 4816 7188 4844 7228
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 6546 7256 6552 7268
rect 6227 7228 6552 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 8036 7256 8064 7355
rect 8202 7352 8208 7404
rect 8260 7352 8266 7404
rect 8297 7395 8355 7401
rect 8297 7361 8309 7395
rect 8343 7361 8355 7395
rect 8297 7355 8355 7361
rect 8312 7324 8340 7355
rect 8570 7352 8576 7404
rect 8628 7352 8634 7404
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 8864 7392 8892 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 11514 7488 11520 7540
rect 11572 7528 11578 7540
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 11572 7500 12265 7528
rect 11572 7488 11578 7500
rect 12253 7497 12265 7500
rect 12299 7497 12311 7531
rect 12253 7491 12311 7497
rect 12345 7531 12403 7537
rect 12345 7497 12357 7531
rect 12391 7528 12403 7531
rect 12710 7528 12716 7540
rect 12391 7500 12716 7528
rect 12391 7497 12403 7500
rect 12345 7491 12403 7497
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 13078 7528 13084 7540
rect 12952 7500 13084 7528
rect 12952 7488 12958 7500
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14424 7500 14473 7528
rect 14424 7488 14430 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 15654 7488 15660 7540
rect 15712 7528 15718 7540
rect 15933 7531 15991 7537
rect 15933 7528 15945 7531
rect 15712 7500 15945 7528
rect 15712 7488 15718 7500
rect 15933 7497 15945 7500
rect 15979 7497 15991 7531
rect 15933 7491 15991 7497
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 17954 7528 17960 7540
rect 16899 7500 17960 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17954 7488 17960 7500
rect 18012 7528 18018 7540
rect 19702 7528 19708 7540
rect 18012 7500 19708 7528
rect 18012 7488 18018 7500
rect 19702 7488 19708 7500
rect 19760 7488 19766 7540
rect 20070 7488 20076 7540
rect 20128 7488 20134 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 22094 7528 22100 7540
rect 20680 7500 21220 7528
rect 20680 7488 20686 7500
rect 8956 7432 9444 7460
rect 8956 7401 8984 7432
rect 8711 7364 8892 7392
rect 8941 7395 8999 7401
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 9217 7355 9275 7361
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8312 7296 9045 7324
rect 9033 7293 9045 7296
rect 9079 7324 9091 7327
rect 9122 7324 9128 7336
rect 9079 7296 9128 7324
rect 9079 7293 9091 7296
rect 9033 7287 9091 7293
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 7116 7228 8064 7256
rect 8849 7259 8907 7265
rect 7116 7197 7144 7228
rect 8849 7225 8861 7259
rect 8895 7256 8907 7259
rect 9232 7256 9260 7355
rect 9416 7333 9444 7432
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 9640 7432 10640 7460
rect 9640 7420 9646 7432
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 10226 7392 10232 7404
rect 10183 7364 10232 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10612 7401 10640 7432
rect 10870 7420 10876 7472
rect 10928 7460 10934 7472
rect 10928 7432 11192 7460
rect 10928 7420 10934 7432
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 11054 7392 11060 7404
rect 11011 7364 11060 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 11164 7401 11192 7432
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 14185 7463 14243 7469
rect 12676 7432 13124 7460
rect 12676 7420 12682 7432
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11238 7392 11244 7404
rect 11195 7364 11244 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11238 7352 11244 7364
rect 11296 7352 11302 7404
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 11974 7392 11980 7404
rect 11931 7364 11980 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 9858 7324 9864 7336
rect 9447 7296 9864 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 9968 7296 10640 7324
rect 9968 7256 9996 7296
rect 8895 7228 9996 7256
rect 8895 7225 8907 7228
rect 8849 7219 8907 7225
rect 10502 7216 10508 7268
rect 10560 7216 10566 7268
rect 10612 7256 10640 7296
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 11422 7256 11428 7268
rect 10612 7228 11428 7256
rect 11422 7216 11428 7228
rect 11480 7256 11486 7268
rect 11900 7256 11928 7355
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12084 7324 12112 7355
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12400 7364 12541 7392
rect 12400 7352 12406 7364
rect 12529 7361 12541 7364
rect 12575 7361 12587 7395
rect 12529 7355 12587 7361
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 13096 7401 13124 7432
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14642 7460 14648 7472
rect 14231 7432 14648 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13596 7364 13829 7392
rect 13596 7352 13602 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 13910 7395 13968 7401
rect 13910 7361 13922 7395
rect 13956 7361 13968 7395
rect 13910 7355 13968 7361
rect 12434 7324 12440 7336
rect 12084 7296 12440 7324
rect 12434 7284 12440 7296
rect 12492 7324 12498 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12492 7296 12725 7324
rect 12492 7284 12498 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 11480 7228 11928 7256
rect 12728 7256 12756 7287
rect 12802 7284 12808 7336
rect 12860 7284 12866 7336
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 13925 7324 13953 7355
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 14056 7364 14105 7392
rect 14056 7352 14062 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 13780 7296 13953 7324
rect 13780 7284 13786 7296
rect 14200 7256 14228 7423
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 18417 7463 18475 7469
rect 18417 7460 18429 7463
rect 15672 7432 18429 7460
rect 14323 7395 14381 7401
rect 14323 7361 14335 7395
rect 14369 7392 14381 7395
rect 14458 7392 14464 7404
rect 14369 7364 14464 7392
rect 14369 7361 14381 7364
rect 14323 7355 14381 7361
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 15672 7401 15700 7432
rect 18417 7429 18429 7432
rect 18463 7429 18475 7463
rect 19886 7460 19892 7472
rect 18417 7423 18475 7429
rect 19444 7432 19892 7460
rect 15657 7395 15715 7401
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15657 7355 15715 7361
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16794 7395 16852 7401
rect 16794 7392 16806 7395
rect 16632 7364 16806 7392
rect 16632 7352 16638 7364
rect 16794 7361 16806 7364
rect 16840 7392 16852 7395
rect 16840 7364 17264 7392
rect 16840 7361 16852 7364
rect 16794 7355 16852 7361
rect 15286 7284 15292 7336
rect 15344 7284 15350 7336
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 12728 7228 14228 7256
rect 15764 7256 15792 7287
rect 16669 7259 16727 7265
rect 16669 7256 16681 7259
rect 15764 7228 16681 7256
rect 11480 7216 11486 7228
rect 16669 7225 16681 7228
rect 16715 7225 16727 7259
rect 17236 7256 17264 7364
rect 17586 7352 17592 7404
rect 17644 7352 17650 7404
rect 17678 7352 17684 7404
rect 17736 7352 17742 7404
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 17954 7352 17960 7404
rect 18012 7352 18018 7404
rect 19444 7401 19472 7432
rect 19886 7420 19892 7432
rect 19944 7420 19950 7472
rect 20898 7460 20904 7472
rect 20364 7432 20904 7460
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7361 19487 7395
rect 19429 7355 19487 7361
rect 17313 7327 17371 7333
rect 17313 7293 17325 7327
rect 17359 7324 17371 7327
rect 18046 7324 18052 7336
rect 17359 7296 18052 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18601 7327 18659 7333
rect 18601 7293 18613 7327
rect 18647 7293 18659 7327
rect 18601 7287 18659 7293
rect 18616 7256 18644 7287
rect 18690 7284 18696 7336
rect 18748 7284 18754 7336
rect 19061 7327 19119 7333
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 19153 7327 19211 7333
rect 19153 7324 19165 7327
rect 19107 7296 19165 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 19153 7293 19165 7296
rect 19199 7293 19211 7327
rect 19352 7324 19380 7355
rect 19702 7352 19708 7404
rect 19760 7352 19766 7404
rect 19518 7324 19524 7336
rect 19352 7296 19524 7324
rect 19153 7287 19211 7293
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 19904 7324 19932 7420
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20364 7401 20392 7432
rect 20898 7420 20904 7432
rect 20956 7420 20962 7472
rect 21192 7469 21220 7500
rect 21284 7500 22100 7528
rect 21284 7469 21312 7500
rect 22094 7488 22100 7500
rect 22152 7488 22158 7540
rect 22278 7488 22284 7540
rect 22336 7528 22342 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 22336 7500 22385 7528
rect 22336 7488 22342 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 22373 7491 22431 7497
rect 22465 7531 22523 7537
rect 22465 7497 22477 7531
rect 22511 7528 22523 7531
rect 22646 7528 22652 7540
rect 22511 7500 22652 7528
rect 22511 7497 22523 7500
rect 22465 7491 22523 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 24210 7488 24216 7540
rect 24268 7528 24274 7540
rect 24581 7531 24639 7537
rect 24581 7528 24593 7531
rect 24268 7500 24593 7528
rect 24268 7488 24274 7500
rect 24581 7497 24593 7500
rect 24627 7497 24639 7531
rect 24581 7491 24639 7497
rect 21177 7463 21235 7469
rect 21177 7429 21189 7463
rect 21223 7429 21235 7463
rect 21177 7423 21235 7429
rect 21269 7463 21327 7469
rect 21269 7429 21281 7463
rect 21315 7429 21327 7463
rect 21269 7423 21327 7429
rect 21542 7420 21548 7472
rect 21600 7460 21606 7472
rect 21910 7460 21916 7472
rect 21600 7432 21916 7460
rect 21600 7420 21606 7432
rect 21910 7420 21916 7432
rect 21968 7460 21974 7472
rect 24670 7460 24676 7472
rect 21968 7432 22140 7460
rect 21968 7420 21974 7432
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20128 7364 20269 7392
rect 20128 7352 20134 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 20625 7395 20683 7401
rect 20625 7361 20637 7395
rect 20671 7361 20683 7395
rect 20625 7355 20683 7361
rect 20640 7324 20668 7355
rect 20990 7352 20996 7404
rect 21048 7392 21054 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 21048 7364 21097 7392
rect 21048 7352 21054 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21450 7352 21456 7404
rect 21508 7352 21514 7404
rect 21818 7352 21824 7404
rect 21876 7392 21882 7404
rect 22112 7401 22140 7432
rect 24320 7432 24676 7460
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21876 7364 22017 7392
rect 21876 7352 21882 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22098 7395 22156 7401
rect 22098 7361 22110 7395
rect 22144 7361 22156 7395
rect 22098 7355 22156 7361
rect 22740 7395 22798 7401
rect 22740 7361 22752 7395
rect 22786 7361 22798 7395
rect 22740 7355 22798 7361
rect 19904 7296 20668 7324
rect 22756 7324 22784 7355
rect 22830 7352 22836 7404
rect 22888 7352 22894 7404
rect 23290 7352 23296 7404
rect 23348 7392 23354 7404
rect 24320 7401 24348 7432
rect 24670 7420 24676 7432
rect 24728 7420 24734 7472
rect 24029 7395 24087 7401
rect 24029 7392 24041 7395
rect 23348 7364 24041 7392
rect 23348 7352 23354 7364
rect 24029 7361 24041 7364
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 23106 7324 23112 7336
rect 22756 7296 23112 7324
rect 23106 7284 23112 7296
rect 23164 7284 23170 7336
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24121 7327 24179 7333
rect 24121 7324 24133 7327
rect 23900 7296 24133 7324
rect 23900 7284 23906 7296
rect 24121 7293 24133 7296
rect 24167 7324 24179 7327
rect 24578 7324 24584 7336
rect 24167 7296 24584 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 29822 7324 29828 7336
rect 24636 7296 29828 7324
rect 24636 7284 24642 7296
rect 29822 7284 29828 7296
rect 29880 7284 29886 7336
rect 20901 7259 20959 7265
rect 20901 7256 20913 7259
rect 17236 7228 17632 7256
rect 18616 7228 20913 7256
rect 16669 7219 16727 7225
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 4816 7160 7113 7188
rect 7101 7157 7113 7160
rect 7147 7157 7159 7191
rect 7101 7151 7159 7157
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 8386 7148 8392 7200
rect 8444 7148 8450 7200
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10962 7188 10968 7200
rect 9916 7160 10968 7188
rect 9916 7148 9922 7160
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 17218 7148 17224 7200
rect 17276 7148 17282 7200
rect 17405 7191 17463 7197
rect 17405 7157 17417 7191
rect 17451 7188 17463 7191
rect 17494 7188 17500 7200
rect 17451 7160 17500 7188
rect 17451 7157 17463 7160
rect 17405 7151 17463 7157
rect 17494 7148 17500 7160
rect 17552 7148 17558 7200
rect 17604 7188 17632 7228
rect 20901 7225 20913 7228
rect 20947 7225 20959 7259
rect 20901 7219 20959 7225
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 17604 7160 19625 7188
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 19613 7151 19671 7157
rect 19702 7148 19708 7200
rect 19760 7188 19766 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 19760 7160 20545 7188
rect 19760 7148 19766 7160
rect 20533 7157 20545 7160
rect 20579 7188 20591 7191
rect 21174 7188 21180 7200
rect 20579 7160 21180 7188
rect 20579 7157 20591 7160
rect 20533 7151 20591 7157
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 1104 7098 29716 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 29716 7098
rect 1104 7024 29716 7046
rect 1670 6993 1676 6996
rect 1660 6987 1676 6993
rect 1660 6953 1672 6987
rect 1660 6947 1676 6953
rect 1670 6944 1676 6947
rect 1728 6944 1734 6996
rect 2958 6944 2964 6996
rect 3016 6984 3022 6996
rect 3145 6987 3203 6993
rect 3145 6984 3157 6987
rect 3016 6956 3157 6984
rect 3016 6944 3022 6956
rect 3145 6953 3157 6956
rect 3191 6953 3203 6987
rect 3145 6947 3203 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 7800 6956 8217 6984
rect 7800 6944 7806 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6984 10195 6987
rect 10226 6984 10232 6996
rect 10183 6956 10232 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 12802 6984 12808 6996
rect 12759 6956 12808 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 15286 6944 15292 6996
rect 15344 6944 15350 6996
rect 17954 6944 17960 6996
rect 18012 6984 18018 6996
rect 18598 6984 18604 6996
rect 18012 6956 18604 6984
rect 18012 6944 18018 6956
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 18877 6987 18935 6993
rect 18877 6984 18889 6987
rect 18748 6956 18889 6984
rect 18748 6944 18754 6956
rect 18877 6953 18889 6956
rect 18923 6953 18935 6987
rect 18877 6947 18935 6953
rect 6822 6876 6828 6928
rect 6880 6916 6886 6928
rect 9766 6916 9772 6928
rect 6880 6888 9772 6916
rect 6880 6876 6886 6888
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 12621 6919 12679 6925
rect 12621 6916 12633 6919
rect 12544 6888 12633 6916
rect 1302 6808 1308 6860
rect 1360 6848 1366 6860
rect 1397 6851 1455 6857
rect 1397 6848 1409 6851
rect 1360 6820 1409 6848
rect 1360 6808 1366 6820
rect 1397 6817 1409 6820
rect 1443 6848 1455 6851
rect 4062 6848 4068 6860
rect 1443 6820 4068 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4614 6848 4620 6860
rect 4571 6820 4620 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8386 6848 8392 6860
rect 8036 6820 8392 6848
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 4706 6780 4712 6792
rect 4479 6752 4712 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 8036 6789 8064 6820
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 12342 6848 12348 6860
rect 10643 6820 12348 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8536 6752 9137 6780
rect 8536 6740 8542 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 2406 6672 2412 6724
rect 2464 6672 2470 6724
rect 4798 6604 4804 6656
rect 4856 6604 4862 6656
rect 9140 6644 9168 6743
rect 9214 6740 9220 6792
rect 9272 6780 9278 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9272 6752 9321 6780
rect 9272 6740 9278 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 10318 6740 10324 6792
rect 10376 6740 10382 6792
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10962 6780 10968 6792
rect 10735 6752 10968 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 12066 6780 12072 6792
rect 11716 6752 12072 6780
rect 10336 6712 10364 6740
rect 11716 6712 11744 6752
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 10336 6684 11744 6712
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 12253 6715 12311 6721
rect 12253 6712 12265 6715
rect 11848 6684 12265 6712
rect 11848 6672 11854 6684
rect 12253 6681 12265 6684
rect 12299 6681 12311 6715
rect 12253 6675 12311 6681
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 12544 6712 12572 6888
rect 12621 6885 12633 6888
rect 12667 6885 12679 6919
rect 12621 6879 12679 6885
rect 13004 6888 13584 6916
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 13004 6857 13032 6888
rect 12989 6851 13047 6857
rect 12989 6848 13001 6851
rect 12768 6820 13001 6848
rect 12768 6808 12774 6820
rect 12989 6817 13001 6820
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13136 6820 13461 6848
rect 13136 6808 13142 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13556 6848 13584 6888
rect 18432 6888 18644 6916
rect 13556 6820 13860 6848
rect 13449 6811 13507 6817
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12676 6752 12909 6780
rect 12676 6740 12682 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13173 6783 13231 6789
rect 13173 6749 13185 6783
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 13188 6712 13216 6743
rect 13262 6740 13268 6792
rect 13320 6780 13326 6792
rect 13357 6783 13415 6789
rect 13357 6780 13369 6783
rect 13320 6752 13369 6780
rect 13320 6740 13326 6752
rect 13357 6749 13369 6752
rect 13403 6749 13415 6783
rect 13464 6780 13492 6811
rect 13832 6789 13860 6820
rect 15010 6808 15016 6860
rect 15068 6848 15074 6860
rect 15068 6820 15700 6848
rect 15068 6808 15074 6820
rect 13633 6783 13691 6789
rect 13633 6780 13645 6783
rect 13464 6752 13645 6780
rect 13357 6743 13415 6749
rect 13633 6749 13645 6752
rect 13679 6749 13691 6783
rect 13633 6743 13691 6749
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6749 13875 6783
rect 13817 6743 13875 6749
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 15286 6712 15292 6724
rect 12544 6684 13216 6712
rect 13280 6684 15292 6712
rect 11698 6644 11704 6656
rect 9140 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 12360 6644 12388 6672
rect 13280 6644 13308 6684
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 15488 6712 15516 6743
rect 15562 6740 15568 6792
rect 15620 6740 15626 6792
rect 15672 6780 15700 6820
rect 15746 6808 15752 6860
rect 15804 6808 15810 6860
rect 16301 6851 16359 6857
rect 16301 6817 16313 6851
rect 16347 6848 16359 6851
rect 16758 6848 16764 6860
rect 16347 6820 16764 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16758 6808 16764 6820
rect 16816 6848 16822 6860
rect 17218 6848 17224 6860
rect 16816 6820 17224 6848
rect 16816 6808 16822 6820
rect 17218 6808 17224 6820
rect 17276 6808 17282 6860
rect 17954 6848 17960 6860
rect 17420 6820 17960 6848
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15672 6752 15853 6780
rect 15841 6749 15853 6752
rect 15887 6780 15899 6783
rect 16114 6780 16120 6792
rect 15887 6752 16120 6780
rect 15887 6749 15899 6752
rect 15841 6743 15899 6749
rect 16114 6740 16120 6752
rect 16172 6740 16178 6792
rect 16206 6740 16212 6792
rect 16264 6740 16270 6792
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6780 17003 6783
rect 17420 6780 17448 6820
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 16991 6752 17448 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 17494 6740 17500 6792
rect 17552 6740 17558 6792
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6780 17831 6783
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17819 6752 18061 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6780 18383 6783
rect 18432 6780 18460 6888
rect 18506 6808 18512 6860
rect 18564 6808 18570 6860
rect 18616 6848 18644 6888
rect 18892 6888 19840 6916
rect 18892 6848 18920 6888
rect 19518 6848 19524 6860
rect 18616 6820 18920 6848
rect 18371 6752 18460 6780
rect 18371 6749 18383 6752
rect 18325 6743 18383 6749
rect 18598 6740 18604 6792
rect 18656 6740 18662 6792
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6780 18843 6783
rect 18892 6780 18920 6820
rect 18984 6820 19524 6848
rect 18984 6789 19012 6820
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 19702 6808 19708 6860
rect 19760 6808 19766 6860
rect 18831 6752 18920 6780
rect 18969 6783 19027 6789
rect 18831 6749 18843 6752
rect 18785 6743 18843 6749
rect 18969 6749 18981 6783
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 19242 6740 19248 6792
rect 19300 6780 19306 6792
rect 19429 6783 19487 6789
rect 19429 6780 19441 6783
rect 19300 6752 19441 6780
rect 19300 6740 19306 6752
rect 19429 6749 19441 6752
rect 19475 6749 19487 6783
rect 19720 6780 19748 6808
rect 19812 6789 19840 6888
rect 20070 6876 20076 6928
rect 20128 6916 20134 6928
rect 20128 6888 21220 6916
rect 20128 6876 20134 6888
rect 19429 6743 19487 6749
rect 19536 6752 19748 6780
rect 19797 6783 19855 6789
rect 16224 6712 16252 6740
rect 15488 6684 16252 6712
rect 16666 6672 16672 6724
rect 16724 6712 16730 6724
rect 16761 6715 16819 6721
rect 16761 6712 16773 6715
rect 16724 6684 16773 6712
rect 16724 6672 16730 6684
rect 16761 6681 16773 6684
rect 16807 6681 16819 6715
rect 17586 6712 17592 6724
rect 16761 6675 16819 6681
rect 16868 6684 17592 6712
rect 12360 6616 13308 6644
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 14090 6644 14096 6656
rect 13771 6616 14096 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15654 6644 15660 6656
rect 15252 6616 15660 6644
rect 15252 6604 15258 6616
rect 15654 6604 15660 6616
rect 15712 6644 15718 6656
rect 16868 6644 16896 6684
rect 17586 6672 17592 6684
rect 17644 6672 17650 6724
rect 19536 6721 19564 6752
rect 19797 6749 19809 6783
rect 19843 6780 19855 6783
rect 19886 6780 19892 6792
rect 19843 6752 19892 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 21192 6789 21220 6888
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 17681 6715 17739 6721
rect 17681 6681 17693 6715
rect 17727 6712 17739 6715
rect 19521 6715 19579 6721
rect 17727 6684 19472 6712
rect 17727 6681 17739 6684
rect 17681 6675 17739 6681
rect 15712 6616 16896 6644
rect 17129 6647 17187 6653
rect 15712 6604 15718 6616
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17218 6644 17224 6656
rect 17175 6616 17224 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17310 6604 17316 6656
rect 17368 6604 17374 6656
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 19334 6644 19340 6656
rect 19291 6616 19340 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19444 6644 19472 6684
rect 19521 6681 19533 6715
rect 19567 6681 19579 6715
rect 19521 6675 19579 6681
rect 19610 6672 19616 6724
rect 19668 6672 19674 6724
rect 19702 6672 19708 6724
rect 19760 6712 19766 6724
rect 23934 6712 23940 6724
rect 19760 6684 23940 6712
rect 19760 6672 19766 6684
rect 23934 6672 23940 6684
rect 23992 6672 23998 6724
rect 20162 6644 20168 6656
rect 19444 6616 20168 6644
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 21082 6604 21088 6656
rect 21140 6604 21146 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 29086 6644 29092 6656
rect 21416 6616 29092 6644
rect 21416 6604 21422 6616
rect 29086 6604 29092 6616
rect 29144 6604 29150 6656
rect 1104 6554 29716 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 29716 6554
rect 1104 6480 29716 6502
rect 2406 6400 2412 6452
rect 2464 6400 2470 6452
rect 8113 6443 8171 6449
rect 8113 6409 8125 6443
rect 8159 6440 8171 6443
rect 8202 6440 8208 6452
rect 8159 6412 8208 6440
rect 8159 6409 8171 6412
rect 8113 6403 8171 6409
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 8478 6440 8484 6452
rect 8312 6412 8484 6440
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 8312 6313 8340 6412
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9180 6412 11928 6440
rect 9180 6400 9186 6412
rect 11900 6384 11928 6412
rect 12618 6400 12624 6452
rect 12676 6400 12682 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 12952 6412 13369 6440
rect 12952 6400 12958 6412
rect 13357 6409 13369 6412
rect 13403 6409 13415 6443
rect 17310 6440 17316 6452
rect 13357 6403 13415 6409
rect 15856 6412 17316 6440
rect 8389 6375 8447 6381
rect 8389 6341 8401 6375
rect 8435 6372 8447 6375
rect 10229 6375 10287 6381
rect 10229 6372 10241 6375
rect 8435 6344 10241 6372
rect 8435 6341 8447 6344
rect 8389 6335 8447 6341
rect 10229 6341 10241 6344
rect 10275 6372 10287 6375
rect 10410 6372 10416 6384
rect 10275 6344 10416 6372
rect 10275 6341 10287 6344
rect 10229 6335 10287 6341
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 11790 6332 11796 6384
rect 11848 6332 11854 6384
rect 11882 6332 11888 6384
rect 11940 6332 11946 6384
rect 11992 6344 15792 6372
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8481 6307 8539 6313
rect 8481 6273 8493 6307
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1719 6208 2774 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2746 6168 2774 6208
rect 6638 6196 6644 6248
rect 6696 6196 6702 6248
rect 8496 6236 8524 6267
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8628 6276 8677 6304
rect 8628 6264 8634 6276
rect 8665 6273 8677 6276
rect 8711 6304 8723 6307
rect 9490 6304 9496 6316
rect 8711 6276 9496 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 9490 6264 9496 6276
rect 9548 6304 9554 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9548 6276 9965 6304
rect 9548 6264 9554 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 9122 6236 9128 6248
rect 6840 6208 9128 6236
rect 6840 6168 6868 6208
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 9968 6236 9996 6267
rect 10134 6264 10140 6316
rect 10192 6264 10198 6316
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6304 10379 6307
rect 11146 6304 11152 6316
rect 10367 6276 11152 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 10962 6236 10968 6248
rect 9968 6208 10968 6236
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 11992 6236 12020 6344
rect 12066 6264 12072 6316
rect 12124 6304 12130 6316
rect 13556 6313 13584 6344
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12124 6276 12449 6304
rect 12124 6264 12130 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6273 13599 6307
rect 13541 6267 13599 6273
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 11112 6208 12265 6236
rect 11112 6196 11118 6208
rect 12253 6205 12265 6208
rect 12299 6205 12311 6239
rect 12452 6236 12480 6267
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 13740 6236 13768 6264
rect 12452 6208 13768 6236
rect 12253 6199 12311 6205
rect 13814 6196 13820 6248
rect 13872 6196 13878 6248
rect 14752 6236 14780 6267
rect 15010 6264 15016 6316
rect 15068 6304 15074 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15068 6276 15301 6304
rect 15068 6264 15074 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 14752 6208 15332 6236
rect 2746 6140 6868 6168
rect 6917 6171 6975 6177
rect 6917 6137 6929 6171
rect 6963 6168 6975 6171
rect 7006 6168 7012 6180
rect 6963 6140 7012 6168
rect 6963 6137 6975 6140
rect 6917 6131 6975 6137
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 15105 6171 15163 6177
rect 15105 6168 15117 6171
rect 8812 6140 15117 6168
rect 8812 6128 8818 6140
rect 15105 6137 15117 6140
rect 15151 6137 15163 6171
rect 15304 6168 15332 6208
rect 15378 6196 15384 6248
rect 15436 6236 15442 6248
rect 15473 6239 15531 6245
rect 15473 6236 15485 6239
rect 15436 6208 15485 6236
rect 15436 6196 15442 6208
rect 15473 6205 15485 6208
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 15562 6196 15568 6248
rect 15620 6196 15626 6248
rect 15764 6236 15792 6344
rect 15856 6313 15884 6412
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 20312 6412 20392 6440
rect 20312 6400 20318 6412
rect 17126 6332 17132 6384
rect 17184 6332 17190 6384
rect 17218 6332 17224 6384
rect 17276 6332 17282 6384
rect 17586 6372 17592 6384
rect 17328 6344 17592 6372
rect 15841 6307 15899 6313
rect 15841 6273 15853 6307
rect 15887 6273 15899 6307
rect 15841 6267 15899 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17328 6304 17356 6344
rect 17586 6332 17592 6344
rect 17644 6332 17650 6384
rect 18230 6332 18236 6384
rect 18288 6372 18294 6384
rect 20364 6381 20392 6412
rect 20732 6412 22385 6440
rect 20349 6375 20407 6381
rect 18288 6344 19564 6372
rect 18288 6332 18294 6344
rect 17083 6276 17356 6304
rect 17405 6307 17463 6313
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17405 6273 17417 6307
rect 17451 6304 17463 6307
rect 19426 6304 19432 6316
rect 17451 6276 19432 6304
rect 17451 6273 17463 6276
rect 17405 6267 17463 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19536 6304 19564 6344
rect 20349 6341 20361 6375
rect 20395 6341 20407 6375
rect 20349 6335 20407 6341
rect 19886 6304 19892 6316
rect 19536 6276 19892 6304
rect 19886 6264 19892 6276
rect 19944 6304 19950 6316
rect 20119 6307 20177 6313
rect 20119 6304 20131 6307
rect 19944 6276 20131 6304
rect 19944 6264 19950 6276
rect 20119 6273 20131 6276
rect 20165 6273 20177 6307
rect 20119 6267 20177 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6273 20315 6307
rect 20257 6267 20315 6273
rect 19702 6236 19708 6248
rect 15764 6208 19708 6236
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 19794 6196 19800 6248
rect 19852 6236 19858 6248
rect 20272 6236 20300 6267
rect 20438 6264 20444 6316
rect 20496 6313 20502 6316
rect 20496 6307 20545 6313
rect 20496 6273 20499 6307
rect 20533 6273 20545 6307
rect 20496 6267 20545 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6304 20683 6307
rect 20732 6304 20760 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 22664 6412 24164 6440
rect 21177 6375 21235 6381
rect 21177 6372 21189 6375
rect 20671 6276 20760 6304
rect 21008 6344 21189 6372
rect 20671 6273 20683 6276
rect 20625 6267 20683 6273
rect 20496 6264 20502 6267
rect 21008 6236 21036 6344
rect 21177 6341 21189 6344
rect 21223 6341 21235 6375
rect 21177 6335 21235 6341
rect 21269 6375 21327 6381
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 21634 6372 21640 6384
rect 21315 6344 21640 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 21634 6332 21640 6344
rect 21692 6332 21698 6384
rect 21080 6307 21138 6313
rect 21080 6273 21092 6307
rect 21126 6304 21138 6307
rect 21126 6276 21220 6304
rect 21126 6273 21138 6276
rect 21080 6267 21138 6273
rect 21192 6248 21220 6276
rect 21450 6264 21456 6316
rect 21508 6264 21514 6316
rect 21542 6264 21548 6316
rect 21600 6264 21606 6316
rect 21818 6264 21824 6316
rect 21876 6264 21882 6316
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 22189 6307 22247 6313
rect 22189 6273 22201 6307
rect 22235 6304 22247 6307
rect 22554 6304 22560 6316
rect 22235 6276 22560 6304
rect 22235 6273 22247 6276
rect 22189 6267 22247 6273
rect 19852 6208 21036 6236
rect 19852 6196 19858 6208
rect 21174 6196 21180 6248
rect 21232 6196 21238 6248
rect 22112 6236 22140 6267
rect 22554 6264 22560 6276
rect 22612 6264 22618 6316
rect 22664 6313 22692 6412
rect 24029 6375 24087 6381
rect 24029 6372 24041 6375
rect 22756 6344 24041 6372
rect 22649 6307 22707 6313
rect 22649 6273 22661 6307
rect 22695 6273 22707 6307
rect 22649 6267 22707 6273
rect 22756 6236 22784 6344
rect 24029 6341 24041 6344
rect 24075 6341 24087 6375
rect 24029 6335 24087 6341
rect 24136 6316 24164 6412
rect 24486 6400 24492 6452
rect 24544 6440 24550 6452
rect 24544 6412 25084 6440
rect 24544 6400 24550 6412
rect 25056 6372 25084 6412
rect 24228 6344 24808 6372
rect 25056 6344 25176 6372
rect 22830 6264 22836 6316
rect 22888 6264 22894 6316
rect 22925 6307 22983 6313
rect 22925 6273 22937 6307
rect 22971 6273 22983 6307
rect 22925 6267 22983 6273
rect 23017 6307 23075 6313
rect 23017 6273 23029 6307
rect 23063 6304 23075 6307
rect 23198 6306 23204 6316
rect 23124 6304 23204 6306
rect 23063 6278 23204 6304
rect 23063 6276 23152 6278
rect 23063 6273 23075 6276
rect 23017 6267 23075 6273
rect 22112 6208 22784 6236
rect 15580 6168 15608 6196
rect 17126 6168 17132 6180
rect 15304 6140 17132 6168
rect 15105 6131 15163 6137
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 20254 6128 20260 6180
rect 20312 6168 20318 6180
rect 21913 6171 21971 6177
rect 21913 6168 21925 6171
rect 20312 6140 21925 6168
rect 20312 6128 20318 6140
rect 21913 6137 21925 6140
rect 21959 6137 21971 6171
rect 21913 6131 21971 6137
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 10284 6072 10517 6100
rect 10284 6060 10290 6072
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 10505 6063 10563 6069
rect 11517 6103 11575 6109
rect 11517 6069 11529 6103
rect 11563 6100 11575 6103
rect 11698 6100 11704 6112
rect 11563 6072 11704 6100
rect 11563 6069 11575 6072
rect 11517 6063 11575 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 11848 6072 14473 6100
rect 11848 6060 11854 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 14918 6060 14924 6112
rect 14976 6060 14982 6112
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 17034 6100 17040 6112
rect 16899 6072 17040 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 17034 6060 17040 6072
rect 17092 6060 17098 6112
rect 18230 6060 18236 6112
rect 18288 6100 18294 6112
rect 19981 6103 20039 6109
rect 19981 6100 19993 6103
rect 18288 6072 19993 6100
rect 18288 6060 18294 6072
rect 19981 6069 19993 6072
rect 20027 6069 20039 6103
rect 19981 6063 20039 6069
rect 20162 6060 20168 6112
rect 20220 6100 20226 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20220 6072 20913 6100
rect 20220 6060 20226 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 22940 6100 22968 6267
rect 23198 6264 23204 6278
rect 23256 6264 23262 6316
rect 23293 6305 23351 6311
rect 23293 6271 23305 6305
rect 23339 6271 23351 6305
rect 23293 6265 23351 6271
rect 23201 6171 23259 6177
rect 23201 6137 23213 6171
rect 23247 6168 23259 6171
rect 23308 6168 23336 6265
rect 23474 6264 23480 6316
rect 23532 6264 23538 6316
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 23750 6304 23756 6316
rect 23707 6276 23756 6304
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 23750 6264 23756 6276
rect 23808 6264 23814 6316
rect 23842 6264 23848 6316
rect 23900 6264 23906 6316
rect 24118 6264 24124 6316
rect 24176 6264 24182 6316
rect 23569 6239 23627 6245
rect 23569 6205 23581 6239
rect 23615 6205 23627 6239
rect 23860 6236 23888 6264
rect 24228 6236 24256 6344
rect 24302 6264 24308 6316
rect 24360 6264 24366 6316
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6273 24455 6307
rect 24397 6267 24455 6273
rect 23860 6208 24256 6236
rect 24412 6236 24440 6267
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 24780 6313 24808 6344
rect 25148 6313 25176 6344
rect 24765 6307 24823 6313
rect 24765 6273 24777 6307
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 25041 6307 25099 6313
rect 25041 6273 25053 6307
rect 25087 6273 25099 6307
rect 25041 6267 25099 6273
rect 25133 6307 25191 6313
rect 25133 6273 25145 6307
rect 25179 6273 25191 6307
rect 25133 6267 25191 6273
rect 25056 6236 25084 6267
rect 29086 6264 29092 6316
rect 29144 6264 29150 6316
rect 24412 6208 25084 6236
rect 23569 6199 23627 6205
rect 23247 6140 23336 6168
rect 23584 6168 23612 6199
rect 23934 6168 23940 6180
rect 23584 6140 23940 6168
rect 23247 6137 23259 6140
rect 23201 6131 23259 6137
rect 23584 6100 23612 6140
rect 23934 6128 23940 6140
rect 23992 6168 23998 6180
rect 24412 6168 24440 6208
rect 29362 6196 29368 6248
rect 29420 6196 29426 6248
rect 23992 6140 24440 6168
rect 23992 6128 23998 6140
rect 24578 6128 24584 6180
rect 24636 6168 24642 6180
rect 24857 6171 24915 6177
rect 24857 6168 24869 6171
rect 24636 6140 24869 6168
rect 24636 6128 24642 6140
rect 24857 6137 24869 6140
rect 24903 6137 24915 6171
rect 24857 6131 24915 6137
rect 22940 6072 23612 6100
rect 24673 6103 24731 6109
rect 20901 6063 20959 6069
rect 24673 6069 24685 6103
rect 24719 6100 24731 6103
rect 24762 6100 24768 6112
rect 24719 6072 24768 6100
rect 24719 6069 24731 6072
rect 24673 6063 24731 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 24946 6060 24952 6112
rect 25004 6100 25010 6112
rect 25317 6103 25375 6109
rect 25317 6100 25329 6103
rect 25004 6072 25329 6100
rect 25004 6060 25010 6072
rect 25317 6069 25329 6072
rect 25363 6069 25375 6103
rect 25317 6063 25375 6069
rect 1104 6010 29716 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 29716 6010
rect 1104 5936 29716 5958
rect 8294 5856 8300 5908
rect 8352 5856 8358 5908
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 11146 5896 11152 5908
rect 10192 5868 11152 5896
rect 10192 5856 10198 5868
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 11514 5856 11520 5908
rect 11572 5856 11578 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13814 5896 13820 5908
rect 13587 5868 13820 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 13964 5868 16129 5896
rect 13964 5856 13970 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16540 5868 16620 5896
rect 16540 5856 16546 5868
rect 8113 5831 8171 5837
rect 8113 5797 8125 5831
rect 8159 5828 8171 5831
rect 8570 5828 8576 5840
rect 8159 5800 8576 5828
rect 8159 5797 8171 5800
rect 8113 5791 8171 5797
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 8665 5831 8723 5837
rect 8665 5797 8677 5831
rect 8711 5828 8723 5831
rect 8941 5831 8999 5837
rect 8941 5828 8953 5831
rect 8711 5800 8953 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 8941 5797 8953 5800
rect 8987 5797 8999 5831
rect 8941 5791 8999 5797
rect 10597 5831 10655 5837
rect 10597 5797 10609 5831
rect 10643 5828 10655 5831
rect 11054 5828 11060 5840
rect 10643 5800 11060 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 14185 5831 14243 5837
rect 14185 5828 14197 5831
rect 11992 5800 14197 5828
rect 3142 5720 3148 5772
rect 3200 5760 3206 5772
rect 5442 5760 5448 5772
rect 3200 5732 5448 5760
rect 3200 5720 3206 5732
rect 5442 5720 5448 5732
rect 5500 5760 5506 5772
rect 7193 5763 7251 5769
rect 7193 5760 7205 5763
rect 5500 5732 7205 5760
rect 5500 5720 5506 5732
rect 7193 5729 7205 5732
rect 7239 5760 7251 5763
rect 7466 5760 7472 5772
rect 7239 5732 7472 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 8754 5720 8760 5772
rect 8812 5720 8818 5772
rect 11606 5760 11612 5772
rect 10060 5732 11612 5760
rect 4154 5652 4160 5704
rect 4212 5652 4218 5704
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7374 5692 7380 5704
rect 7147 5664 7380 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7374 5652 7380 5664
rect 7432 5692 7438 5704
rect 8018 5692 8024 5704
rect 7432 5664 8024 5692
rect 7432 5652 7438 5664
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8478 5652 8484 5704
rect 8536 5652 8542 5704
rect 8938 5652 8944 5704
rect 8996 5692 9002 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8996 5664 9137 5692
rect 8996 5652 9002 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9214 5652 9220 5704
rect 9272 5692 9278 5704
rect 10060 5701 10088 5732
rect 11606 5720 11612 5732
rect 11664 5720 11670 5772
rect 11992 5760 12020 5800
rect 14185 5797 14197 5800
rect 14231 5797 14243 5831
rect 14185 5791 14243 5797
rect 15470 5788 15476 5840
rect 15528 5828 15534 5840
rect 15528 5800 16528 5828
rect 15528 5788 15534 5800
rect 16500 5769 16528 5800
rect 16592 5769 16620 5868
rect 16666 5856 16672 5908
rect 16724 5896 16730 5908
rect 17310 5896 17316 5908
rect 16724 5868 17316 5896
rect 16724 5856 16730 5868
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 18506 5896 18512 5908
rect 17460 5868 18512 5896
rect 17460 5856 17466 5868
rect 18506 5856 18512 5868
rect 18564 5896 18570 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 18564 5868 18889 5896
rect 18564 5856 18570 5868
rect 18877 5865 18889 5868
rect 18923 5865 18935 5899
rect 18877 5859 18935 5865
rect 19242 5856 19248 5908
rect 19300 5896 19306 5908
rect 19794 5896 19800 5908
rect 19300 5868 19800 5896
rect 19300 5856 19306 5868
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 19904 5868 22094 5896
rect 18598 5828 18604 5840
rect 16684 5800 18604 5828
rect 16485 5763 16543 5769
rect 11900 5732 12020 5760
rect 14568 5732 16436 5760
rect 9493 5695 9551 5701
rect 9272 5664 9444 5692
rect 9272 5652 9278 5664
rect 4430 5584 4436 5636
rect 4488 5584 4494 5636
rect 8846 5584 8852 5636
rect 8904 5624 8910 5636
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8904 5596 9321 5624
rect 8904 5584 8910 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 9416 5624 9444 5664
rect 9493 5661 9505 5695
rect 9539 5692 9551 5695
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9539 5664 10057 5692
rect 9539 5661 9551 5664
rect 9493 5655 9551 5661
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10318 5692 10324 5704
rect 10045 5655 10103 5661
rect 10152 5664 10324 5692
rect 9582 5624 9588 5636
rect 9416 5596 9588 5624
rect 9309 5587 9367 5593
rect 9582 5584 9588 5596
rect 9640 5624 9646 5636
rect 10152 5624 10180 5664
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10410 5652 10416 5704
rect 10468 5692 10474 5704
rect 10873 5695 10931 5701
rect 10873 5692 10885 5695
rect 10468 5664 10885 5692
rect 10468 5652 10474 5664
rect 10873 5661 10885 5664
rect 10919 5661 10931 5695
rect 10873 5655 10931 5661
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11698 5652 11704 5704
rect 11756 5652 11762 5704
rect 11900 5701 11928 5732
rect 11885 5695 11943 5701
rect 11885 5661 11897 5695
rect 11931 5661 11943 5695
rect 11885 5655 11943 5661
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13078 5701 13084 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12676 5664 12909 5692
rect 12676 5652 12682 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 13045 5695 13084 5701
rect 13045 5661 13057 5695
rect 13045 5655 13084 5661
rect 13078 5652 13084 5655
rect 13136 5652 13142 5704
rect 13446 5701 13452 5704
rect 13403 5695 13452 5701
rect 13403 5661 13415 5695
rect 13449 5661 13452 5695
rect 13403 5655 13452 5661
rect 13446 5652 13452 5655
rect 13504 5652 13510 5704
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 14568 5701 14596 5732
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 13872 5664 14381 5692
rect 13872 5652 13878 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 14642 5652 14648 5704
rect 14700 5652 14706 5704
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 16301 5695 16359 5701
rect 16301 5692 16313 5695
rect 15804 5664 16313 5692
rect 15804 5652 15810 5664
rect 16301 5661 16313 5664
rect 16347 5661 16359 5695
rect 16301 5655 16359 5661
rect 9640 5596 10180 5624
rect 10229 5627 10287 5633
rect 9640 5584 9646 5596
rect 10229 5593 10241 5627
rect 10275 5593 10287 5627
rect 10229 5587 10287 5593
rect 5902 5516 5908 5568
rect 5960 5516 5966 5568
rect 6638 5516 6644 5568
rect 6696 5516 6702 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10244 5556 10272 5587
rect 13170 5584 13176 5636
rect 13228 5584 13234 5636
rect 13262 5584 13268 5636
rect 13320 5624 13326 5636
rect 15654 5624 15660 5636
rect 13320 5596 15660 5624
rect 13320 5584 13326 5596
rect 15654 5584 15660 5596
rect 15712 5584 15718 5636
rect 10192 5528 10272 5556
rect 10192 5516 10198 5528
rect 10686 5516 10692 5568
rect 10744 5516 10750 5568
rect 16316 5556 16344 5655
rect 16408 5624 16436 5732
rect 16485 5729 16497 5763
rect 16531 5729 16543 5763
rect 16485 5723 16543 5729
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5729 16635 5763
rect 16577 5723 16635 5729
rect 16684 5701 16712 5800
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 16776 5732 17877 5760
rect 16669 5695 16727 5701
rect 16669 5661 16681 5695
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 16776 5624 16804 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 19904 5760 19932 5868
rect 21085 5831 21143 5837
rect 21085 5797 21097 5831
rect 21131 5828 21143 5831
rect 21542 5828 21548 5840
rect 21131 5800 21548 5828
rect 21131 5797 21143 5800
rect 21085 5791 21143 5797
rect 21542 5788 21548 5800
rect 21600 5788 21606 5840
rect 22066 5828 22094 5868
rect 22554 5856 22560 5908
rect 22612 5856 22618 5908
rect 29638 5828 29644 5840
rect 22066 5800 29644 5828
rect 29638 5788 29644 5800
rect 29696 5788 29702 5840
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 17865 5723 17923 5729
rect 17972 5732 19932 5760
rect 20456 5732 21649 5760
rect 16850 5652 16856 5704
rect 16908 5652 16914 5704
rect 17218 5652 17224 5704
rect 17276 5652 17282 5704
rect 17402 5652 17408 5704
rect 17460 5652 17466 5704
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5692 17647 5695
rect 17678 5692 17684 5704
rect 17635 5664 17684 5692
rect 17635 5661 17647 5664
rect 17589 5655 17647 5661
rect 17678 5652 17684 5664
rect 17736 5652 17742 5704
rect 16408 5596 16804 5624
rect 17494 5584 17500 5636
rect 17552 5584 17558 5636
rect 17972 5624 18000 5732
rect 20456 5704 20484 5732
rect 21637 5729 21649 5732
rect 21683 5760 21695 5763
rect 21818 5760 21824 5772
rect 21683 5732 21824 5760
rect 21683 5729 21695 5732
rect 21637 5723 21695 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 23750 5760 23756 5772
rect 22756 5732 23756 5760
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 17604 5596 18000 5624
rect 17604 5556 17632 5596
rect 16316 5528 17632 5556
rect 17773 5559 17831 5565
rect 17773 5525 17785 5559
rect 17819 5556 17831 5559
rect 18064 5556 18092 5655
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 18371 5664 18429 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5692 19027 5695
rect 19058 5692 19064 5704
rect 19015 5664 19064 5692
rect 19015 5661 19027 5664
rect 18969 5655 19027 5661
rect 17819 5528 18092 5556
rect 18616 5556 18644 5655
rect 18708 5624 18736 5655
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 19576 5664 19717 5692
rect 19576 5652 19582 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5692 20131 5695
rect 20438 5692 20444 5704
rect 20119 5664 20444 5692
rect 20119 5661 20131 5664
rect 20073 5655 20131 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 20901 5695 20959 5701
rect 20901 5661 20913 5695
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 19242 5624 19248 5636
rect 18708 5596 19248 5624
rect 19242 5584 19248 5596
rect 19300 5584 19306 5636
rect 19996 5624 20024 5652
rect 20640 5624 20668 5655
rect 19996 5596 20668 5624
rect 20916 5624 20944 5655
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21140 5664 21189 5692
rect 21140 5652 21146 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 22756 5701 22784 5732
rect 23750 5720 23756 5732
rect 23808 5720 23814 5772
rect 21729 5695 21787 5701
rect 21729 5692 21741 5695
rect 21416 5664 21741 5692
rect 21416 5652 21422 5664
rect 21729 5661 21741 5664
rect 21775 5661 21787 5695
rect 21729 5655 21787 5661
rect 22741 5695 22799 5701
rect 22741 5661 22753 5695
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 22922 5652 22928 5704
rect 22980 5692 22986 5704
rect 23842 5692 23848 5704
rect 22980 5664 23848 5692
rect 22980 5652 22986 5664
rect 23842 5652 23848 5664
rect 23900 5692 23906 5704
rect 23900 5664 24532 5692
rect 23900 5652 23906 5664
rect 21376 5624 21404 5652
rect 20916 5596 21404 5624
rect 21450 5584 21456 5636
rect 21508 5624 21514 5636
rect 24504 5624 24532 5664
rect 24578 5652 24584 5704
rect 24636 5652 24642 5704
rect 24762 5652 24768 5704
rect 24820 5652 24826 5704
rect 24946 5652 24952 5704
rect 25004 5652 25010 5704
rect 24673 5627 24731 5633
rect 24673 5624 24685 5627
rect 21508 5596 24440 5624
rect 24504 5596 24685 5624
rect 21508 5584 21514 5596
rect 19702 5556 19708 5568
rect 18616 5528 19708 5556
rect 17819 5525 17831 5528
rect 17773 5519 17831 5525
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 20070 5516 20076 5568
rect 20128 5556 20134 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 20128 5528 20269 5556
rect 20128 5516 20134 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 20990 5556 20996 5568
rect 20763 5528 20996 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 20990 5516 20996 5528
rect 21048 5556 21054 5568
rect 21266 5556 21272 5568
rect 21048 5528 21272 5556
rect 21048 5516 21054 5528
rect 21266 5516 21272 5528
rect 21324 5516 21330 5568
rect 21361 5559 21419 5565
rect 21361 5525 21373 5559
rect 21407 5556 21419 5559
rect 21634 5556 21640 5568
rect 21407 5528 21640 5556
rect 21407 5525 21419 5528
rect 21361 5519 21419 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 24412 5565 24440 5596
rect 24673 5593 24685 5596
rect 24719 5593 24731 5627
rect 24673 5587 24731 5593
rect 24397 5559 24455 5565
rect 24397 5525 24409 5559
rect 24443 5525 24455 5559
rect 24397 5519 24455 5525
rect 1104 5466 29716 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 29716 5466
rect 1104 5392 29716 5414
rect 4430 5312 4436 5364
rect 4488 5352 4494 5364
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 4488 5324 4721 5352
rect 4488 5312 4494 5324
rect 4709 5321 4721 5324
rect 4755 5321 4767 5355
rect 4709 5315 4767 5321
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 5077 5355 5135 5361
rect 5077 5352 5089 5355
rect 4856 5324 5089 5352
rect 4856 5312 4862 5324
rect 5077 5321 5089 5324
rect 5123 5321 5135 5355
rect 5077 5315 5135 5321
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5592 5324 5641 5352
rect 5592 5312 5598 5324
rect 5629 5321 5641 5324
rect 5675 5321 5687 5355
rect 5629 5315 5687 5321
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 8076 5324 8125 5352
rect 8076 5312 8082 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8113 5315 8171 5321
rect 8478 5312 8484 5364
rect 8536 5352 8542 5364
rect 8757 5355 8815 5361
rect 8757 5352 8769 5355
rect 8536 5324 8769 5352
rect 8536 5312 8542 5324
rect 8757 5321 8769 5324
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 10008 5324 10057 5352
rect 10008 5312 10014 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10045 5315 10103 5321
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11974 5352 11980 5364
rect 11563 5324 11980 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 13814 5352 13820 5364
rect 12759 5324 13820 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 14090 5312 14096 5364
rect 14148 5312 14154 5364
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14700 5324 14933 5352
rect 14700 5312 14706 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 16482 5312 16488 5364
rect 16540 5312 16546 5364
rect 16850 5312 16856 5364
rect 16908 5312 16914 5364
rect 18141 5355 18199 5361
rect 18141 5321 18153 5355
rect 18187 5352 18199 5355
rect 20162 5352 20168 5364
rect 18187 5324 20168 5352
rect 18187 5321 18199 5324
rect 18141 5315 18199 5321
rect 20162 5312 20168 5324
rect 20220 5312 20226 5364
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 22097 5355 22155 5361
rect 22097 5352 22109 5355
rect 20487 5324 22109 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 22097 5321 22109 5324
rect 22143 5321 22155 5355
rect 22097 5315 22155 5321
rect 22186 5312 22192 5364
rect 22244 5312 22250 5364
rect 23934 5312 23940 5364
rect 23992 5312 23998 5364
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 5902 5284 5908 5296
rect 5215 5256 5908 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 5902 5244 5908 5256
rect 5960 5244 5966 5296
rect 6638 5244 6644 5296
rect 6696 5244 6702 5296
rect 8297 5287 8355 5293
rect 8297 5284 8309 5287
rect 7866 5256 8309 5284
rect 8297 5253 8309 5256
rect 8343 5253 8355 5287
rect 8297 5247 8355 5253
rect 8570 5244 8576 5296
rect 8628 5284 8634 5296
rect 10413 5287 10471 5293
rect 8628 5256 9352 5284
rect 8628 5244 8634 5256
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 900 5188 1501 5216
rect 900 5176 906 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4212 5188 5580 5216
rect 4212 5176 4218 5188
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5148 5411 5151
rect 5442 5148 5448 5160
rect 5399 5120 5448 5148
rect 5399 5117 5411 5120
rect 5353 5111 5411 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5552 5148 5580 5188
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5684 5188 5733 5216
rect 5684 5176 5690 5188
rect 5721 5185 5733 5188
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5185 8447 5219
rect 8389 5179 8447 5185
rect 6362 5148 6368 5160
rect 5552 5120 6368 5148
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 8404 5148 8432 5179
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5216 9091 5219
rect 9214 5216 9220 5228
rect 9079 5188 9220 5216
rect 9079 5185 9091 5188
rect 9033 5179 9091 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9324 5225 9352 5256
rect 10413 5253 10425 5287
rect 10459 5284 10471 5287
rect 10873 5287 10931 5293
rect 10873 5284 10885 5287
rect 10459 5256 10885 5284
rect 10459 5253 10471 5256
rect 10413 5247 10471 5253
rect 10873 5253 10885 5256
rect 10919 5253 10931 5287
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 10873 5247 10931 5253
rect 11716 5256 12940 5284
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10686 5216 10692 5228
rect 10551 5188 10692 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11054 5176 11060 5228
rect 11112 5176 11118 5228
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 11333 5219 11391 5225
rect 11333 5185 11345 5219
rect 11379 5216 11391 5219
rect 11606 5216 11612 5228
rect 11379 5188 11612 5216
rect 11379 5185 11391 5188
rect 11333 5179 11391 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11716 5225 11744 5256
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11793 5222 11851 5225
rect 11793 5219 11928 5222
rect 11793 5185 11805 5219
rect 11839 5216 11928 5219
rect 11974 5216 11980 5228
rect 11839 5194 11980 5216
rect 11839 5185 11851 5194
rect 11900 5188 11980 5194
rect 11793 5179 11851 5185
rect 6472 5120 8432 5148
rect 8956 5148 8984 5176
rect 11716 5148 11744 5179
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 12912 5225 12940 5256
rect 13372 5256 14197 5284
rect 12897 5219 12955 5225
rect 12897 5185 12909 5219
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 12989 5219 13047 5225
rect 12989 5185 13001 5219
rect 13035 5185 13047 5219
rect 12989 5179 13047 5185
rect 8956 5120 11744 5148
rect 11992 5148 12020 5176
rect 13004 5148 13032 5179
rect 13078 5176 13084 5228
rect 13136 5176 13142 5228
rect 13262 5176 13268 5228
rect 13320 5176 13326 5228
rect 13372 5225 13400 5256
rect 14185 5253 14197 5256
rect 14231 5253 14243 5287
rect 14185 5247 14243 5253
rect 14553 5287 14611 5293
rect 14553 5253 14565 5287
rect 14599 5284 14611 5287
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 14599 5256 17785 5284
rect 14599 5253 14611 5256
rect 14553 5247 14611 5253
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 18598 5244 18604 5296
rect 18656 5244 18662 5296
rect 22204 5284 22232 5312
rect 22373 5287 22431 5293
rect 22373 5284 22385 5287
rect 18892 5256 20300 5284
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 13538 5176 13544 5228
rect 13596 5176 13602 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13872 5188 13921 5216
rect 13872 5176 13878 5188
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 14366 5176 14372 5228
rect 14424 5176 14430 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5216 14703 5219
rect 14826 5216 14832 5228
rect 14691 5188 14832 5216
rect 14691 5185 14703 5188
rect 14645 5179 14703 5185
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 15102 5176 15108 5228
rect 15160 5176 15166 5228
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15243 5188 15424 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 13446 5148 13452 5160
rect 11992 5120 13452 5148
rect 5626 5040 5632 5092
rect 5684 5080 5690 5092
rect 6472 5080 6500 5120
rect 5684 5052 6500 5080
rect 8404 5080 8432 5120
rect 13446 5108 13452 5120
rect 13504 5148 13510 5160
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 13504 5120 13645 5148
rect 13504 5108 13510 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5148 13783 5151
rect 13998 5148 14004 5160
rect 13771 5120 14004 5148
rect 13771 5117 13783 5120
rect 13725 5111 13783 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 15010 5108 15016 5160
rect 15068 5148 15074 5160
rect 15396 5148 15424 5188
rect 15470 5176 15476 5228
rect 15528 5176 15534 5228
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15620 5188 15945 5216
rect 15620 5176 15626 5188
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16114 5176 16120 5228
rect 16172 5176 16178 5228
rect 16206 5176 16212 5228
rect 16264 5176 16270 5228
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16316 5148 16344 5179
rect 16666 5176 16672 5228
rect 16724 5176 16730 5228
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16816 5188 16865 5216
rect 16816 5176 16822 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17218 5216 17224 5228
rect 17175 5188 17224 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17310 5176 17316 5228
rect 17368 5176 17374 5228
rect 17402 5176 17408 5228
rect 17460 5176 17466 5228
rect 17497 5219 17555 5225
rect 17497 5185 17509 5219
rect 17543 5216 17555 5219
rect 17586 5216 17592 5228
rect 17543 5188 17592 5216
rect 17543 5185 17555 5188
rect 17497 5179 17555 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17696 5188 17969 5216
rect 17420 5148 17448 5176
rect 15068 5120 17448 5148
rect 15068 5108 15074 5120
rect 9030 5080 9036 5092
rect 8404 5052 9036 5080
rect 5684 5040 5690 5052
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9217 5083 9275 5089
rect 9217 5080 9229 5083
rect 9180 5052 9229 5080
rect 9180 5040 9186 5052
rect 9217 5049 9229 5052
rect 9263 5049 9275 5083
rect 9217 5043 9275 5049
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 11296 5052 12434 5080
rect 11296 5040 11302 5052
rect 1578 4972 1584 5024
rect 1636 4972 1642 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11940 4984 11989 5012
rect 11940 4972 11946 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 12406 5012 12434 5052
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 15378 5080 15384 5092
rect 13136 5052 15384 5080
rect 13136 5040 13142 5052
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 16114 5040 16120 5092
rect 16172 5080 16178 5092
rect 17218 5080 17224 5092
rect 16172 5052 17224 5080
rect 16172 5040 16178 5052
rect 17218 5040 17224 5052
rect 17276 5040 17282 5092
rect 17696 5089 17724 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18506 5216 18512 5228
rect 18279 5188 18512 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18892 5225 18920 5256
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 18877 5219 18935 5225
rect 18877 5185 18889 5219
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 18800 5148 18828 5179
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 19153 5219 19211 5225
rect 19153 5216 19165 5219
rect 19024 5188 19165 5216
rect 19024 5176 19030 5188
rect 19153 5185 19165 5188
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19334 5176 19340 5228
rect 19392 5216 19398 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 19392 5188 19441 5216
rect 19392 5176 19398 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 20070 5176 20076 5228
rect 20128 5176 20134 5228
rect 20272 5225 20300 5256
rect 21192 5256 22385 5284
rect 21192 5225 21220 5256
rect 22373 5253 22385 5256
rect 22419 5253 22431 5287
rect 22373 5247 22431 5253
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 20533 5219 20591 5225
rect 20533 5185 20545 5219
rect 20579 5216 20591 5219
rect 20901 5219 20959 5225
rect 20901 5216 20913 5219
rect 20579 5188 20913 5216
rect 20579 5185 20591 5188
rect 20533 5179 20591 5185
rect 20901 5185 20913 5188
rect 20947 5185 20959 5219
rect 20901 5179 20959 5185
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 21177 5219 21235 5225
rect 21177 5185 21189 5219
rect 21223 5185 21235 5219
rect 21177 5179 21235 5185
rect 19245 5151 19303 5157
rect 19245 5148 19257 5151
rect 18800 5120 19257 5148
rect 19245 5117 19257 5120
rect 19291 5117 19303 5151
rect 21100 5148 21128 5179
rect 21266 5176 21272 5228
rect 21324 5216 21330 5228
rect 22278 5225 22284 5228
rect 21453 5219 21511 5225
rect 21453 5216 21465 5219
rect 21324 5188 21465 5216
rect 21324 5176 21330 5188
rect 21453 5185 21465 5188
rect 21499 5185 21511 5219
rect 22235 5219 22284 5225
rect 22235 5216 22247 5219
rect 21453 5179 21511 5185
rect 22066 5188 22247 5216
rect 22066 5148 22094 5188
rect 22235 5185 22247 5188
rect 22281 5185 22284 5219
rect 22235 5179 22284 5185
rect 22278 5176 22284 5179
rect 22336 5176 22342 5228
rect 22462 5176 22468 5228
rect 22520 5176 22526 5228
rect 22646 5176 22652 5228
rect 22704 5176 22710 5228
rect 22738 5176 22744 5228
rect 22796 5176 22802 5228
rect 23842 5176 23848 5228
rect 23900 5216 23906 5228
rect 24029 5219 24087 5225
rect 24029 5216 24041 5219
rect 23900 5188 24041 5216
rect 23900 5176 23906 5188
rect 24029 5185 24041 5188
rect 24075 5185 24087 5219
rect 24029 5179 24087 5185
rect 29270 5176 29276 5228
rect 29328 5176 29334 5228
rect 21100 5120 22094 5148
rect 19245 5111 19303 5117
rect 17681 5083 17739 5089
rect 17681 5049 17693 5083
rect 17727 5049 17739 5083
rect 18966 5080 18972 5092
rect 17681 5043 17739 5049
rect 18708 5052 18972 5080
rect 17034 5012 17040 5024
rect 12406 4984 17040 5012
rect 11977 4975 12035 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 18708 5012 18736 5052
rect 18966 5040 18972 5052
rect 19024 5040 19030 5092
rect 19058 5040 19064 5092
rect 19116 5040 19122 5092
rect 29089 5083 29147 5089
rect 29089 5080 29101 5083
rect 19168 5052 29101 5080
rect 17184 4984 18736 5012
rect 17184 4972 17190 4984
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19168 5012 19196 5052
rect 29089 5049 29101 5052
rect 29135 5049 29147 5083
rect 29089 5043 29147 5049
rect 18840 4984 19196 5012
rect 18840 4972 18846 4984
rect 21082 4972 21088 5024
rect 21140 5012 21146 5024
rect 21358 5012 21364 5024
rect 21140 4984 21364 5012
rect 21140 4972 21146 4984
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 1104 4922 29716 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 29716 4922
rect 1104 4848 29716 4870
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 13078 4808 13084 4820
rect 8904 4780 13084 4808
rect 8904 4768 8910 4780
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13817 4811 13875 4817
rect 13464 4780 13768 4808
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 10042 4740 10048 4752
rect 1636 4712 10048 4740
rect 1636 4700 1642 4712
rect 10042 4700 10048 4712
rect 10100 4700 10106 4752
rect 10134 4700 10140 4752
rect 10192 4740 10198 4752
rect 11977 4743 12035 4749
rect 10192 4712 11928 4740
rect 10192 4700 10198 4712
rect 11900 4672 11928 4712
rect 11977 4709 11989 4743
rect 12023 4740 12035 4743
rect 12066 4740 12072 4752
rect 12023 4712 12072 4740
rect 12023 4709 12035 4712
rect 11977 4703 12035 4709
rect 12066 4700 12072 4712
rect 12124 4700 12130 4752
rect 13464 4672 13492 4780
rect 13740 4740 13768 4780
rect 13817 4777 13829 4811
rect 13863 4808 13875 4811
rect 14366 4808 14372 4820
rect 13863 4780 14372 4808
rect 13863 4777 13875 4780
rect 13817 4771 13875 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14826 4768 14832 4820
rect 14884 4768 14890 4820
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 14976 4780 15301 4808
rect 14976 4768 14982 4780
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15289 4771 15347 4777
rect 15562 4768 15568 4820
rect 15620 4808 15626 4820
rect 16574 4808 16580 4820
rect 15620 4780 16580 4808
rect 15620 4768 15626 4780
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 16853 4811 16911 4817
rect 16853 4777 16865 4811
rect 16899 4808 16911 4811
rect 17402 4808 17408 4820
rect 16899 4780 17408 4808
rect 16899 4777 16911 4780
rect 16853 4771 16911 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 18506 4768 18512 4820
rect 18564 4768 18570 4820
rect 22373 4811 22431 4817
rect 22373 4777 22385 4811
rect 22419 4808 22431 4811
rect 22738 4808 22744 4820
rect 22419 4780 22744 4808
rect 22419 4777 22431 4780
rect 22373 4771 22431 4777
rect 22738 4768 22744 4780
rect 22796 4768 22802 4820
rect 23937 4811 23995 4817
rect 23937 4777 23949 4811
rect 23983 4808 23995 4811
rect 24118 4808 24124 4820
rect 23983 4780 24124 4808
rect 23983 4777 23995 4780
rect 23937 4771 23995 4777
rect 14936 4740 14964 4768
rect 13740 4712 14964 4740
rect 16592 4740 16620 4768
rect 17126 4740 17132 4752
rect 16592 4712 17132 4740
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 17310 4700 17316 4752
rect 17368 4740 17374 4752
rect 18969 4743 19027 4749
rect 18969 4740 18981 4743
rect 17368 4712 18981 4740
rect 17368 4700 17374 4712
rect 18969 4709 18981 4712
rect 19015 4740 19027 4743
rect 19426 4740 19432 4752
rect 19015 4712 19432 4740
rect 19015 4709 19027 4712
rect 18969 4703 19027 4709
rect 19426 4700 19432 4712
rect 19484 4700 19490 4752
rect 22281 4743 22339 4749
rect 22281 4709 22293 4743
rect 22327 4709 22339 4743
rect 22281 4703 22339 4709
rect 11900 4644 13492 4672
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 11532 4536 11560 4567
rect 11698 4564 11704 4616
rect 11756 4564 11762 4616
rect 11882 4564 11888 4616
rect 11940 4604 11946 4616
rect 12618 4604 12624 4616
rect 11940 4576 12624 4604
rect 11940 4564 11946 4576
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12710 4564 12716 4616
rect 12768 4564 12774 4616
rect 13262 4564 13268 4616
rect 13320 4564 13326 4616
rect 13464 4613 13492 4644
rect 13538 4632 13544 4684
rect 13596 4672 13602 4684
rect 19242 4672 19248 4684
rect 13596 4644 13676 4672
rect 13596 4632 13602 4644
rect 13648 4613 13676 4644
rect 18800 4644 19248 4672
rect 13449 4607 13507 4613
rect 13449 4573 13461 4607
rect 13495 4573 13507 4607
rect 13449 4567 13507 4573
rect 13633 4607 13691 4613
rect 13633 4573 13645 4607
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 14734 4564 14740 4616
rect 14792 4604 14798 4616
rect 15013 4607 15071 4613
rect 15013 4604 15025 4607
rect 14792 4576 15025 4604
rect 14792 4564 14798 4576
rect 15013 4573 15025 4576
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 11974 4536 11980 4548
rect 11532 4508 11980 4536
rect 11974 4496 11980 4508
rect 12032 4536 12038 4548
rect 12250 4536 12256 4548
rect 12032 4508 12256 4536
rect 12032 4496 12038 4508
rect 12250 4496 12256 4508
rect 12308 4536 12314 4548
rect 12805 4539 12863 4545
rect 12805 4536 12817 4539
rect 12308 4508 12817 4536
rect 12308 4496 12314 4508
rect 12805 4505 12817 4508
rect 12851 4536 12863 4539
rect 13541 4539 13599 4545
rect 13541 4536 13553 4539
rect 12851 4508 13553 4536
rect 12851 4505 12863 4508
rect 12805 4499 12863 4505
rect 13541 4505 13553 4508
rect 13587 4505 13599 4539
rect 15028 4536 15056 4567
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15470 4604 15476 4616
rect 15427 4576 15476 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 16666 4564 16672 4616
rect 16724 4604 16730 4616
rect 16761 4607 16819 4613
rect 16761 4604 16773 4607
rect 16724 4576 16773 4604
rect 16724 4564 16730 4576
rect 16761 4573 16773 4576
rect 16807 4604 16819 4607
rect 16850 4604 16856 4616
rect 16807 4576 16856 4604
rect 16807 4573 16819 4576
rect 16761 4567 16819 4573
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 18800 4613 18828 4644
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 22296 4672 22324 4703
rect 22462 4700 22468 4752
rect 22520 4700 22526 4752
rect 22646 4700 22652 4752
rect 22704 4740 22710 4752
rect 22925 4743 22983 4749
rect 22925 4740 22937 4743
rect 22704 4712 22937 4740
rect 22704 4700 22710 4712
rect 22925 4709 22937 4712
rect 22971 4709 22983 4743
rect 22925 4703 22983 4709
rect 23385 4675 23443 4681
rect 21968 4644 22094 4672
rect 22296 4644 22876 4672
rect 21968 4632 21974 4644
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4573 18751 4607
rect 18693 4567 18751 4573
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 17678 4536 17684 4548
rect 15028 4508 17684 4536
rect 13541 4499 13599 4505
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11517 4471 11575 4477
rect 11517 4468 11529 4471
rect 11112 4440 11529 4468
rect 11112 4428 11118 4440
rect 11517 4437 11529 4440
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 11606 4428 11612 4480
rect 11664 4468 11670 4480
rect 17310 4468 17316 4480
rect 11664 4440 17316 4468
rect 11664 4428 11670 4440
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 18708 4468 18736 4567
rect 19058 4564 19064 4616
rect 19116 4564 19122 4616
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 20346 4604 20352 4616
rect 19484 4576 20352 4604
rect 19484 4564 19490 4576
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 22066 4604 22094 4644
rect 22848 4616 22876 4644
rect 23385 4641 23397 4675
rect 23431 4672 23443 4675
rect 23952 4672 23980 4771
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 23431 4644 23980 4672
rect 23431 4641 23443 4644
rect 23385 4635 23443 4641
rect 22679 4607 22737 4613
rect 22679 4604 22691 4607
rect 22066 4576 22691 4604
rect 22679 4573 22691 4576
rect 22725 4573 22737 4607
rect 22679 4567 22737 4573
rect 22830 4564 22836 4616
rect 22888 4564 22894 4616
rect 23106 4564 23112 4616
rect 23164 4613 23170 4616
rect 23164 4607 23197 4613
rect 23185 4573 23197 4607
rect 23164 4567 23197 4573
rect 23293 4607 23351 4613
rect 23293 4573 23305 4607
rect 23339 4604 23351 4607
rect 23474 4604 23480 4616
rect 23339 4576 23480 4604
rect 23339 4573 23351 4576
rect 23293 4567 23351 4573
rect 23164 4564 23170 4567
rect 23474 4564 23480 4576
rect 23532 4564 23538 4616
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 21174 4536 21180 4548
rect 19306 4508 21180 4536
rect 19306 4468 19334 4508
rect 21174 4496 21180 4508
rect 21232 4496 21238 4548
rect 18708 4440 19334 4468
rect 20438 4428 20444 4480
rect 20496 4428 20502 4480
rect 23198 4428 23204 4480
rect 23256 4468 23262 4480
rect 23584 4468 23612 4567
rect 23658 4564 23664 4616
rect 23716 4604 23722 4616
rect 24029 4607 24087 4613
rect 24029 4604 24041 4607
rect 23716 4576 24041 4604
rect 23716 4564 23722 4576
rect 24029 4573 24041 4576
rect 24075 4604 24087 4607
rect 24118 4604 24124 4616
rect 24075 4576 24124 4604
rect 24075 4573 24087 4576
rect 24029 4567 24087 4573
rect 24118 4564 24124 4576
rect 24176 4564 24182 4616
rect 24489 4607 24547 4613
rect 24489 4573 24501 4607
rect 24535 4604 24547 4607
rect 25314 4604 25320 4616
rect 24535 4576 25320 4604
rect 24535 4573 24547 4576
rect 24489 4567 24547 4573
rect 25314 4564 25320 4576
rect 25372 4564 25378 4616
rect 23256 4440 23612 4468
rect 23256 4428 23262 4440
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 24486 4428 24492 4480
rect 24544 4468 24550 4480
rect 24581 4471 24639 4477
rect 24581 4468 24593 4471
rect 24544 4440 24593 4468
rect 24544 4428 24550 4440
rect 24581 4437 24593 4440
rect 24627 4437 24639 4471
rect 24581 4431 24639 4437
rect 1104 4378 29716 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 29716 4378
rect 1104 4304 29716 4326
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11882 4264 11888 4276
rect 10735 4236 11888 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 9950 4156 9956 4208
rect 10008 4156 10014 4208
rect 10962 4156 10968 4208
rect 11020 4196 11026 4208
rect 11164 4205 11192 4236
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 12176 4236 12480 4264
rect 11149 4199 11207 4205
rect 11020 4168 11100 4196
rect 11020 4156 11026 4168
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 6420 4100 8953 4128
rect 6420 4088 6426 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 11072 4128 11100 4168
rect 11149 4165 11161 4199
rect 11195 4165 11207 4199
rect 11149 4159 11207 4165
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 11701 4199 11759 4205
rect 11701 4196 11713 4199
rect 11296 4168 11713 4196
rect 11296 4156 11302 4168
rect 11701 4165 11713 4168
rect 11747 4165 11759 4199
rect 11701 4159 11759 4165
rect 11072 4100 11192 4128
rect 8941 4091 8999 4097
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 11164 4060 11192 4100
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12176 4137 12204 4236
rect 12250 4156 12256 4208
rect 12308 4156 12314 4208
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 11848 4100 12173 4128
rect 11848 4088 11854 4100
rect 12161 4097 12173 4100
rect 12207 4097 12219 4131
rect 12268 4128 12296 4156
rect 12345 4131 12403 4137
rect 12345 4128 12357 4131
rect 12268 4100 12357 4128
rect 12161 4091 12219 4097
rect 12345 4097 12357 4100
rect 12391 4097 12403 4131
rect 12345 4091 12403 4097
rect 12253 4063 12311 4069
rect 12253 4060 12265 4063
rect 9263 4032 10824 4060
rect 11164 4032 12265 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 10796 3924 10824 4032
rect 12253 4029 12265 4032
rect 12299 4029 12311 4063
rect 12452 4060 12480 4236
rect 12710 4224 12716 4276
rect 12768 4224 12774 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 15105 4267 15163 4273
rect 15105 4264 15117 4267
rect 13320 4236 15117 4264
rect 13320 4224 13326 4236
rect 15105 4233 15117 4236
rect 15151 4264 15163 4267
rect 15470 4264 15476 4276
rect 15151 4236 15476 4264
rect 15151 4233 15163 4236
rect 15105 4227 15163 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 17276 4236 17785 4264
rect 17276 4224 17282 4236
rect 17773 4233 17785 4236
rect 17819 4264 17831 4267
rect 19058 4264 19064 4276
rect 17819 4236 19064 4264
rect 17819 4233 17831 4236
rect 17773 4227 17831 4233
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 19153 4267 19211 4273
rect 19153 4233 19165 4267
rect 19199 4264 19211 4267
rect 19242 4264 19248 4276
rect 19199 4236 19248 4264
rect 19199 4233 19211 4236
rect 19153 4227 19211 4233
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 20346 4224 20352 4276
rect 20404 4264 20410 4276
rect 25314 4264 25320 4276
rect 20404 4236 25320 4264
rect 20404 4224 20410 4236
rect 25314 4224 25320 4236
rect 25372 4224 25378 4276
rect 12529 4199 12587 4205
rect 12529 4165 12541 4199
rect 12575 4196 12587 4199
rect 12618 4196 12624 4208
rect 12575 4168 12624 4196
rect 12575 4165 12587 4168
rect 12529 4159 12587 4165
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 12805 4199 12863 4205
rect 12805 4165 12817 4199
rect 12851 4196 12863 4199
rect 12851 4168 13400 4196
rect 12851 4165 12863 4168
rect 12805 4159 12863 4165
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13170 4128 13176 4140
rect 12943 4100 13176 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13372 4137 13400 4168
rect 13814 4156 13820 4208
rect 13872 4196 13878 4208
rect 14550 4196 14556 4208
rect 13872 4168 14556 4196
rect 13872 4156 13878 4168
rect 14550 4156 14556 4168
rect 14608 4196 14614 4208
rect 14737 4199 14795 4205
rect 14737 4196 14749 4199
rect 14608 4168 14749 4196
rect 14608 4156 14614 4168
rect 14737 4165 14749 4168
rect 14783 4196 14795 4199
rect 14783 4168 15148 4196
rect 14783 4165 14795 4168
rect 14737 4159 14795 4165
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13446 4128 13452 4140
rect 13403 4100 13452 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13446 4088 13452 4100
rect 13504 4128 13510 4140
rect 14826 4128 14832 4140
rect 13504 4100 14832 4128
rect 13504 4088 13510 4100
rect 14826 4088 14832 4100
rect 14884 4128 14890 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14884 4100 15025 4128
rect 14884 4088 14890 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 12452 4032 13277 4060
rect 12253 4023 12311 4029
rect 13265 4029 13277 4032
rect 13311 4060 13323 4063
rect 13630 4060 13636 4072
rect 13311 4032 13636 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 14369 4063 14427 4069
rect 14369 4029 14381 4063
rect 14415 4060 14427 4063
rect 15120 4060 15148 4168
rect 16316 4168 16896 4196
rect 16316 4137 16344 4168
rect 16868 4137 16896 4168
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 16531 4100 16681 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16669 4097 16681 4100
rect 16715 4097 16727 4131
rect 16669 4091 16727 4097
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 17236 4128 17264 4224
rect 18064 4168 18276 4196
rect 16899 4100 17264 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 16390 4060 16396 4072
rect 14415 4032 15056 4060
rect 15120 4032 16396 4060
rect 14415 4029 14427 4032
rect 14369 4023 14427 4029
rect 11333 3995 11391 4001
rect 11333 3961 11345 3995
rect 11379 3992 11391 3995
rect 12069 3995 12127 4001
rect 11379 3964 11744 3992
rect 11379 3961 11391 3964
rect 11333 3955 11391 3961
rect 11716 3933 11744 3964
rect 12069 3961 12081 3995
rect 12115 3961 12127 3995
rect 12069 3955 12127 3961
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 10796 3896 11529 3924
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3893 11759 3927
rect 12084 3924 12112 3955
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 14384 3992 14412 4023
rect 13228 3964 14412 3992
rect 13228 3952 13234 3964
rect 14642 3952 14648 4004
rect 14700 3992 14706 4004
rect 14921 3995 14979 4001
rect 14921 3992 14933 3995
rect 14700 3964 14933 3992
rect 14700 3952 14706 3964
rect 14921 3961 14933 3964
rect 14967 3961 14979 3995
rect 15028 3992 15056 4032
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16684 4060 16712 4091
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 17644 4100 17693 4128
rect 17644 4088 17650 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 17957 4131 18015 4137
rect 17957 4097 17969 4131
rect 18003 4128 18015 4131
rect 18064 4128 18092 4168
rect 18248 4140 18276 4168
rect 20438 4156 20444 4208
rect 20496 4156 20502 4208
rect 23750 4156 23756 4208
rect 23808 4156 23814 4208
rect 24486 4156 24492 4208
rect 24544 4156 24550 4208
rect 18003 4100 18092 4128
rect 18003 4097 18015 4100
rect 17957 4091 18015 4097
rect 18138 4088 18144 4140
rect 18196 4088 18202 4140
rect 18230 4088 18236 4140
rect 18288 4128 18294 4140
rect 19061 4131 19119 4137
rect 19061 4128 19073 4131
rect 18288 4100 19073 4128
rect 18288 4088 18294 4100
rect 19061 4097 19073 4100
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19429 4063 19487 4069
rect 16684 4032 18092 4060
rect 17954 3992 17960 4004
rect 15028 3964 17960 3992
rect 14921 3955 14979 3961
rect 17954 3952 17960 3964
rect 18012 3952 18018 4004
rect 18064 3936 18092 4032
rect 19429 4029 19441 4063
rect 19475 4029 19487 4063
rect 19429 4023 19487 4029
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12084 3896 13093 3924
rect 11701 3887 11759 3893
rect 13081 3893 13093 3896
rect 13127 3924 13139 3927
rect 13354 3924 13360 3936
rect 13127 3896 13360 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 14734 3884 14740 3936
rect 14792 3884 14798 3936
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16574 3924 16580 3936
rect 16439 3896 16580 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16666 3884 16672 3936
rect 16724 3884 16730 3936
rect 18046 3884 18052 3936
rect 18104 3884 18110 3936
rect 19444 3924 19472 4023
rect 19702 4020 19708 4072
rect 19760 4020 19766 4072
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 23477 4063 23535 4069
rect 23477 4060 23489 4063
rect 23348 4032 23489 4060
rect 23348 4020 23354 4032
rect 23477 4029 23489 4032
rect 23523 4029 23535 4063
rect 23477 4023 23535 4029
rect 20714 3924 20720 3936
rect 19444 3896 20720 3924
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 21082 3884 21088 3936
rect 21140 3924 21146 3936
rect 21177 3927 21235 3933
rect 21177 3924 21189 3927
rect 21140 3896 21189 3924
rect 21140 3884 21146 3896
rect 21177 3893 21189 3896
rect 21223 3924 21235 3927
rect 22554 3924 22560 3936
rect 21223 3896 22560 3924
rect 21223 3893 21235 3896
rect 21177 3887 21235 3893
rect 22554 3884 22560 3896
rect 22612 3884 22618 3936
rect 22646 3884 22652 3936
rect 22704 3924 22710 3936
rect 22922 3924 22928 3936
rect 22704 3896 22928 3924
rect 22704 3884 22710 3896
rect 22922 3884 22928 3896
rect 22980 3924 22986 3936
rect 23382 3924 23388 3936
rect 22980 3896 23388 3924
rect 22980 3884 22986 3896
rect 23382 3884 23388 3896
rect 23440 3884 23446 3936
rect 23492 3924 23520 4023
rect 24118 4020 24124 4072
rect 24176 4060 24182 4072
rect 25225 4063 25283 4069
rect 25225 4060 25237 4063
rect 24176 4032 25237 4060
rect 24176 4020 24182 4032
rect 25225 4029 25237 4032
rect 25271 4029 25283 4063
rect 25225 4023 25283 4029
rect 25038 3924 25044 3936
rect 23492 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 1104 3834 29716 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 29716 3834
rect 1104 3760 29716 3782
rect 9950 3680 9956 3732
rect 10008 3680 10014 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 11054 3720 11060 3732
rect 10735 3692 11060 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 12710 3680 12716 3732
rect 12768 3680 12774 3732
rect 13262 3680 13268 3732
rect 13320 3720 13326 3732
rect 13449 3723 13507 3729
rect 13449 3720 13461 3723
rect 13320 3692 13461 3720
rect 13320 3680 13326 3692
rect 13449 3689 13461 3692
rect 13495 3689 13507 3723
rect 13449 3683 13507 3689
rect 13630 3680 13636 3732
rect 13688 3680 13694 3732
rect 16574 3680 16580 3732
rect 16632 3680 16638 3732
rect 17954 3680 17960 3732
rect 18012 3680 18018 3732
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 18693 3723 18751 3729
rect 18693 3720 18705 3723
rect 18104 3692 18705 3720
rect 18104 3680 18110 3692
rect 18693 3689 18705 3692
rect 18739 3689 18751 3723
rect 18693 3683 18751 3689
rect 19797 3723 19855 3729
rect 19797 3689 19809 3723
rect 19843 3720 19855 3723
rect 20257 3723 20315 3729
rect 20257 3720 20269 3723
rect 19843 3692 20269 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 20257 3689 20269 3692
rect 20303 3689 20315 3723
rect 20257 3683 20315 3689
rect 20824 3692 22722 3720
rect 10321 3655 10379 3661
rect 10321 3621 10333 3655
rect 10367 3652 10379 3655
rect 10962 3652 10968 3664
rect 10367 3624 10968 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 10962 3612 10968 3624
rect 11020 3612 11026 3664
rect 16209 3655 16267 3661
rect 16209 3621 16221 3655
rect 16255 3652 16267 3655
rect 16666 3652 16672 3664
rect 16255 3624 16672 3652
rect 16255 3621 16267 3624
rect 16209 3615 16267 3621
rect 16666 3612 16672 3624
rect 16724 3612 16730 3664
rect 16761 3655 16819 3661
rect 16761 3621 16773 3655
rect 16807 3652 16819 3655
rect 17862 3652 17868 3664
rect 16807 3624 17868 3652
rect 16807 3621 16819 3624
rect 16761 3615 16819 3621
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 18414 3612 18420 3664
rect 18472 3612 18478 3664
rect 18524 3624 19564 3652
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11296 3556 12572 3584
rect 11296 3544 11302 3556
rect 842 3476 848 3528
rect 900 3516 906 3528
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 900 3488 1501 3516
rect 900 3476 906 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9582 3516 9588 3528
rect 9088 3488 9588 3516
rect 9088 3476 9094 3488
rect 9582 3476 9588 3488
rect 9640 3516 9646 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 9640 3488 9873 3516
rect 9640 3476 9646 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3448 10747 3451
rect 11146 3448 11152 3460
rect 10735 3420 11152 3448
rect 10735 3417 10747 3420
rect 10689 3411 10747 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11241 3451 11299 3457
rect 11241 3417 11253 3451
rect 11287 3417 11299 3451
rect 11241 3411 11299 3417
rect 1578 3340 1584 3392
rect 1636 3340 1642 3392
rect 10873 3383 10931 3389
rect 10873 3349 10885 3383
rect 10919 3380 10931 3383
rect 11256 3380 11284 3411
rect 11974 3408 11980 3460
rect 12032 3408 12038 3460
rect 10919 3352 11284 3380
rect 12544 3380 12572 3556
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 14332 3556 14381 3584
rect 14332 3544 14338 3556
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 14642 3544 14648 3596
rect 14700 3544 14706 3596
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 18524 3584 18552 3624
rect 19334 3584 19340 3596
rect 15344 3556 18552 3584
rect 15344 3544 15350 3556
rect 19306 3544 19340 3584
rect 19392 3584 19398 3596
rect 19429 3587 19487 3593
rect 19429 3584 19441 3587
rect 19392 3556 19441 3584
rect 19392 3544 19398 3556
rect 19429 3553 19441 3556
rect 19475 3553 19487 3587
rect 19429 3547 19487 3553
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 13078 3516 13084 3528
rect 13035 3488 13084 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13446 3516 13452 3528
rect 13219 3488 13452 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3516 17739 3519
rect 18230 3516 18236 3528
rect 17727 3488 18236 3516
rect 17727 3485 17739 3488
rect 17681 3479 17739 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 19306 3516 19334 3544
rect 18340 3488 19334 3516
rect 19536 3516 19564 3624
rect 19702 3612 19708 3664
rect 19760 3652 19766 3664
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 19760 3624 19993 3652
rect 19760 3612 19766 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 20824 3652 20852 3692
rect 19981 3615 20039 3621
rect 20088 3624 20852 3652
rect 20088 3516 20116 3624
rect 22278 3612 22284 3664
rect 22336 3652 22342 3664
rect 22462 3652 22468 3664
rect 22336 3624 22468 3652
rect 22336 3612 22342 3624
rect 22462 3612 22468 3624
rect 22520 3612 22526 3664
rect 22554 3612 22560 3664
rect 22612 3612 22618 3664
rect 22694 3652 22722 3692
rect 23106 3680 23112 3732
rect 23164 3680 23170 3732
rect 23293 3723 23351 3729
rect 23293 3689 23305 3723
rect 23339 3720 23351 3723
rect 23382 3720 23388 3732
rect 23339 3692 23388 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 23382 3680 23388 3692
rect 23440 3720 23446 3732
rect 23658 3720 23664 3732
rect 23440 3692 23664 3720
rect 23440 3680 23446 3692
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 29089 3655 29147 3661
rect 29089 3652 29101 3655
rect 22694 3624 29101 3652
rect 29089 3621 29101 3624
rect 29135 3621 29147 3655
rect 29089 3615 29147 3621
rect 21082 3584 21088 3596
rect 20456 3556 21088 3584
rect 20456 3525 20484 3556
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 23382 3584 23388 3596
rect 22796 3556 23388 3584
rect 22796 3544 22802 3556
rect 23382 3544 23388 3556
rect 23440 3584 23446 3596
rect 23845 3587 23903 3593
rect 23845 3584 23857 3587
rect 23440 3556 23857 3584
rect 23440 3544 23446 3556
rect 19536 3488 20116 3516
rect 20441 3519 20499 3525
rect 13357 3451 13415 3457
rect 13357 3417 13369 3451
rect 13403 3448 13415 3451
rect 13601 3451 13659 3457
rect 13601 3448 13613 3451
rect 13403 3420 13613 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 13601 3417 13613 3420
rect 13647 3417 13659 3451
rect 13601 3411 13659 3417
rect 13814 3408 13820 3460
rect 13872 3408 13878 3460
rect 15378 3408 15384 3460
rect 15436 3408 15442 3460
rect 16850 3448 16856 3460
rect 16132 3420 16856 3448
rect 13832 3380 13860 3408
rect 16132 3392 16160 3420
rect 16850 3408 16856 3420
rect 16908 3448 16914 3460
rect 17405 3451 17463 3457
rect 17405 3448 17417 3451
rect 16908 3420 17417 3448
rect 16908 3408 16914 3420
rect 17405 3417 17417 3420
rect 17451 3417 17463 3451
rect 17773 3451 17831 3457
rect 17405 3411 17463 3417
rect 17512 3420 17724 3448
rect 12544 3352 13860 3380
rect 10919 3349 10931 3352
rect 10873 3343 10931 3349
rect 16114 3340 16120 3392
rect 16172 3340 16178 3392
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16577 3383 16635 3389
rect 16577 3380 16589 3383
rect 16448 3352 16589 3380
rect 16448 3340 16454 3352
rect 16577 3349 16589 3352
rect 16623 3380 16635 3383
rect 17512 3380 17540 3420
rect 16623 3352 17540 3380
rect 16623 3349 16635 3352
rect 16577 3343 16635 3349
rect 17586 3340 17592 3392
rect 17644 3340 17650 3392
rect 17696 3380 17724 3420
rect 17773 3417 17785 3451
rect 17819 3448 17831 3451
rect 18049 3451 18107 3457
rect 18049 3448 18061 3451
rect 17819 3420 18061 3448
rect 17819 3417 17831 3420
rect 17773 3411 17831 3417
rect 18049 3417 18061 3420
rect 18095 3448 18107 3451
rect 18138 3448 18144 3460
rect 18095 3420 18144 3448
rect 18095 3417 18107 3420
rect 18049 3411 18107 3417
rect 18138 3408 18144 3420
rect 18196 3448 18202 3460
rect 18340 3448 18368 3488
rect 20441 3485 20453 3519
rect 20487 3485 20499 3519
rect 20441 3479 20499 3485
rect 20714 3476 20720 3528
rect 20772 3476 20778 3528
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 23492 3525 23520 3556
rect 23845 3553 23857 3556
rect 23891 3553 23903 3587
rect 23845 3547 23903 3553
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 22520 3488 23213 3516
rect 22520 3476 22526 3488
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 23750 3476 23756 3528
rect 23808 3476 23814 3528
rect 23937 3519 23995 3525
rect 23937 3485 23949 3519
rect 23983 3516 23995 3519
rect 24118 3516 24124 3528
rect 23983 3488 24124 3516
rect 23983 3485 23995 3488
rect 23937 3479 23995 3485
rect 18196 3420 18368 3448
rect 18509 3451 18567 3457
rect 18196 3408 18202 3420
rect 18509 3417 18521 3451
rect 18555 3448 18567 3451
rect 19797 3451 19855 3457
rect 19797 3448 19809 3451
rect 18555 3420 19809 3448
rect 18555 3417 18567 3420
rect 18509 3411 18567 3417
rect 19797 3417 19809 3420
rect 19843 3448 19855 3451
rect 20346 3448 20352 3460
rect 19843 3420 20352 3448
rect 19843 3417 19855 3420
rect 19797 3411 19855 3417
rect 18524 3380 18552 3411
rect 20346 3408 20352 3420
rect 20404 3408 20410 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 20993 3451 21051 3457
rect 20680 3420 20944 3448
rect 20680 3408 20686 3420
rect 17696 3352 18552 3380
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 18709 3383 18767 3389
rect 18709 3380 18721 3383
rect 18656 3352 18721 3380
rect 18656 3340 18662 3352
rect 18709 3349 18721 3352
rect 18755 3349 18767 3383
rect 18709 3343 18767 3349
rect 18877 3383 18935 3389
rect 18877 3349 18889 3383
rect 18923 3380 18935 3383
rect 19702 3380 19708 3392
rect 18923 3352 19708 3380
rect 18923 3349 18935 3352
rect 18877 3343 18935 3349
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 20916 3380 20944 3420
rect 20993 3417 21005 3451
rect 21039 3448 21051 3451
rect 21266 3448 21272 3460
rect 21039 3420 21272 3448
rect 21039 3417 21051 3420
rect 20993 3411 21051 3417
rect 21266 3408 21272 3420
rect 21324 3408 21330 3460
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23569 3451 23627 3457
rect 23569 3448 23581 3451
rect 22291 3420 23581 3448
rect 22291 3380 22319 3420
rect 23569 3417 23581 3420
rect 23615 3417 23627 3451
rect 23569 3411 23627 3417
rect 20916 3352 22319 3380
rect 22462 3340 22468 3392
rect 22520 3380 22526 3392
rect 22741 3383 22799 3389
rect 22741 3380 22753 3383
rect 22520 3352 22753 3380
rect 22520 3340 22526 3352
rect 22741 3349 22753 3352
rect 22787 3349 22799 3383
rect 22741 3343 22799 3349
rect 22830 3340 22836 3392
rect 22888 3340 22894 3392
rect 22925 3383 22983 3389
rect 22925 3349 22937 3383
rect 22971 3380 22983 3383
rect 23474 3380 23480 3392
rect 22971 3352 23480 3380
rect 22971 3349 22983 3352
rect 22925 3343 22983 3349
rect 23474 3340 23480 3352
rect 23532 3380 23538 3392
rect 23952 3380 23980 3479
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 29270 3408 29276 3460
rect 29328 3408 29334 3460
rect 23532 3352 23980 3380
rect 23532 3340 23538 3352
rect 1104 3290 29716 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 29716 3290
rect 1104 3216 29716 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 1949 3179 2007 3185
rect 1949 3176 1961 3179
rect 1912 3148 1961 3176
rect 1912 3136 1918 3148
rect 1949 3145 1961 3148
rect 1995 3145 2007 3179
rect 1949 3139 2007 3145
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11793 3179 11851 3185
rect 11793 3176 11805 3179
rect 11388 3148 11805 3176
rect 11388 3136 11394 3148
rect 11793 3145 11805 3148
rect 11839 3145 11851 3179
rect 11793 3139 11851 3145
rect 11974 3136 11980 3188
rect 12032 3176 12038 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 12032 3148 12081 3176
rect 12032 3136 12038 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 12069 3139 12127 3145
rect 12158 3136 12164 3188
rect 12216 3176 12222 3188
rect 14274 3176 14280 3188
rect 12216 3148 14280 3176
rect 12216 3136 12222 3148
rect 11698 3108 11704 3120
rect 1872 3080 2774 3108
rect 1872 3049 1900 3080
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3040 1639 3043
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1627 3012 1869 3040
rect 1627 3009 1639 3012
rect 1581 3003 1639 3009
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 2148 2972 2176 3003
rect 716 2944 2176 2972
rect 2746 2972 2774 3080
rect 9646 3080 11704 3108
rect 9646 3052 9674 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 13060 3108 13088 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 14792 3148 15332 3176
rect 14792 3136 14798 3148
rect 13004 3080 13088 3108
rect 9582 3000 9588 3052
rect 9640 3012 9674 3052
rect 11885 3043 11943 3049
rect 11885 3040 11897 3043
rect 11808 3012 11897 3040
rect 9640 3000 9646 3012
rect 11606 2972 11612 2984
rect 2746 2944 11612 2972
rect 716 2932 722 2944
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 842 2864 848 2916
rect 900 2904 906 2916
rect 1673 2907 1731 2913
rect 1673 2904 1685 2907
rect 900 2876 1685 2904
rect 900 2864 906 2876
rect 1673 2873 1685 2876
rect 1719 2873 1731 2907
rect 11514 2904 11520 2916
rect 1673 2867 1731 2873
rect 2746 2876 11520 2904
rect 1578 2796 1584 2848
rect 1636 2836 1642 2848
rect 2746 2836 2774 2876
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 1636 2808 2774 2836
rect 11808 2836 11836 3012
rect 11885 3009 11897 3012
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3038 12035 3043
rect 12066 3038 12072 3052
rect 12023 3010 12072 3038
rect 12023 3009 12035 3010
rect 11977 3003 12035 3009
rect 12066 3000 12072 3010
rect 12124 3000 12130 3052
rect 13004 3049 13032 3080
rect 13262 3068 13268 3120
rect 13320 3068 13326 3120
rect 14921 3111 14979 3117
rect 14921 3108 14933 3111
rect 14490 3080 14933 3108
rect 14921 3077 14933 3080
rect 14967 3077 14979 3111
rect 15304 3108 15332 3148
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 15436 3148 15485 3176
rect 15436 3136 15442 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 18432 3148 20208 3176
rect 15933 3111 15991 3117
rect 15933 3108 15945 3111
rect 15304 3080 15945 3108
rect 14921 3071 14979 3077
rect 15933 3077 15945 3080
rect 15979 3077 15991 3111
rect 15933 3071 15991 3077
rect 16114 3068 16120 3120
rect 16172 3068 16178 3120
rect 16301 3111 16359 3117
rect 16301 3077 16313 3111
rect 16347 3108 16359 3111
rect 16666 3108 16672 3120
rect 16347 3080 16672 3108
rect 16347 3077 16359 3080
rect 16301 3071 16359 3077
rect 16666 3068 16672 3080
rect 16724 3068 16730 3120
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 18141 3111 18199 3117
rect 18141 3108 18153 3111
rect 17920 3080 18153 3108
rect 17920 3068 17926 3080
rect 18141 3077 18153 3080
rect 18187 3077 18199 3111
rect 18141 3071 18199 3077
rect 12989 3043 13047 3049
rect 12989 3009 13001 3043
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 15059 3012 15393 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15381 3009 15393 3012
rect 15427 3040 15439 3043
rect 16482 3040 16488 3052
rect 15427 3012 16488 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 12084 2972 12112 3000
rect 15028 2972 15056 3003
rect 16482 3000 16488 3012
rect 16540 3000 16546 3052
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 18432 3049 18460 3148
rect 19334 3068 19340 3120
rect 19392 3068 19398 3120
rect 19702 3068 19708 3120
rect 19760 3108 19766 3120
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 19760 3080 19993 3108
rect 19760 3068 19766 3080
rect 19981 3077 19993 3080
rect 20027 3077 20039 3111
rect 20180 3108 20208 3148
rect 21266 3136 21272 3188
rect 21324 3136 21330 3188
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3176 21971 3179
rect 22002 3176 22008 3188
rect 21959 3148 22008 3176
rect 21959 3145 21971 3148
rect 21913 3139 21971 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22922 3136 22928 3188
rect 22980 3176 22986 3188
rect 23750 3176 23756 3188
rect 22980 3148 23756 3176
rect 22980 3136 22986 3148
rect 20714 3108 20720 3120
rect 20180 3080 20720 3108
rect 19981 3071 20039 3077
rect 20272 3049 20300 3080
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 21085 3111 21143 3117
rect 21085 3077 21097 3111
rect 21131 3108 21143 3111
rect 22649 3111 22707 3117
rect 22649 3108 22661 3111
rect 21131 3080 22661 3108
rect 21131 3077 21143 3080
rect 21085 3071 21143 3077
rect 22649 3077 22661 3080
rect 22695 3077 22707 3111
rect 22649 3071 22707 3077
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3009 20315 3043
rect 22005 3043 22063 3049
rect 22005 3040 22017 3043
rect 20257 3003 20315 3009
rect 20548 3012 22017 3040
rect 12084 2944 15056 2972
rect 16669 2975 16727 2981
rect 16669 2941 16681 2975
rect 16715 2972 16727 2975
rect 17586 2972 17592 2984
rect 16715 2944 17592 2972
rect 16715 2941 16727 2944
rect 16669 2935 16727 2941
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18196 2944 18521 2972
rect 18196 2932 18202 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 19426 2932 19432 2984
rect 19484 2972 19490 2984
rect 20548 2972 20576 3012
rect 22005 3009 22017 3012
rect 22051 3009 22063 3043
rect 22005 3003 22063 3009
rect 22554 3000 22560 3052
rect 22612 3000 22618 3052
rect 22738 3000 22744 3052
rect 22796 3000 22802 3052
rect 23032 3049 23060 3148
rect 23750 3136 23756 3148
rect 23808 3176 23814 3188
rect 25041 3179 25099 3185
rect 25041 3176 25053 3179
rect 23808 3148 25053 3176
rect 23808 3136 23814 3148
rect 25041 3145 25053 3148
rect 25087 3145 25099 3179
rect 25041 3139 25099 3145
rect 23474 3108 23480 3120
rect 23216 3080 23480 3108
rect 22833 3043 22891 3049
rect 22833 3009 22845 3043
rect 22879 3009 22891 3043
rect 22833 3003 22891 3009
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3009 23075 3043
rect 23017 3003 23075 3009
rect 19484 2944 20576 2972
rect 19484 2932 19490 2944
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 20717 2975 20775 2981
rect 20717 2972 20729 2975
rect 20680 2944 20729 2972
rect 20680 2932 20686 2944
rect 20717 2941 20729 2944
rect 20763 2941 20775 2975
rect 22848 2972 22876 3003
rect 23216 2972 23244 3080
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 25225 3111 25283 3117
rect 25225 3108 25237 3111
rect 24794 3080 25237 3108
rect 25225 3077 25237 3080
rect 25271 3077 25283 3111
rect 25225 3071 25283 3077
rect 28718 3068 28724 3120
rect 28776 3068 28782 3120
rect 23290 3000 23296 3052
rect 23348 3000 23354 3052
rect 25314 3000 25320 3052
rect 25372 3000 25378 3052
rect 28905 3043 28963 3049
rect 28905 3009 28917 3043
rect 28951 3040 28963 3043
rect 28994 3040 29000 3052
rect 28951 3012 29000 3040
rect 28951 3009 28963 3012
rect 28905 3003 28963 3009
rect 28994 3000 29000 3012
rect 29052 3000 29058 3052
rect 29273 3043 29331 3049
rect 29273 3009 29285 3043
rect 29319 3040 29331 3043
rect 29362 3040 29368 3052
rect 29319 3012 29368 3040
rect 29319 3009 29331 3012
rect 29273 3003 29331 3009
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 22848 2944 23244 2972
rect 20717 2935 20775 2941
rect 23566 2932 23572 2984
rect 23624 2932 23630 2984
rect 22002 2904 22008 2916
rect 14292 2876 14872 2904
rect 11882 2836 11888 2848
rect 11808 2808 11888 2836
rect 1636 2796 1642 2808
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 14292 2836 14320 2876
rect 12032 2808 14320 2836
rect 12032 2796 12038 2808
rect 14734 2796 14740 2848
rect 14792 2796 14798 2848
rect 14844 2836 14872 2876
rect 20180 2876 22008 2904
rect 20180 2836 20208 2876
rect 22002 2864 22008 2876
rect 22060 2864 22066 2916
rect 22922 2904 22928 2916
rect 22480 2876 22928 2904
rect 14844 2808 20208 2836
rect 20346 2796 20352 2848
rect 20404 2836 20410 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 20404 2808 21097 2836
rect 20404 2796 20410 2808
rect 21085 2805 21097 2808
rect 21131 2836 21143 2839
rect 22480 2836 22508 2876
rect 22922 2864 22928 2876
rect 22980 2864 22986 2916
rect 29086 2864 29092 2916
rect 29144 2864 29150 2916
rect 21131 2808 22508 2836
rect 23201 2839 23259 2845
rect 21131 2805 21143 2808
rect 21085 2799 21143 2805
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23382 2836 23388 2848
rect 23247 2808 23388 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 1104 2746 29716 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 29716 2746
rect 1104 2672 29716 2694
rect 8202 2632 8208 2644
rect 2332 2604 8208 2632
rect 2332 2505 2360 2604
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 8297 2635 8355 2641
rect 8297 2601 8309 2635
rect 8343 2632 8355 2635
rect 8662 2632 8668 2644
rect 8343 2604 8668 2632
rect 8343 2601 8355 2604
rect 8297 2595 8355 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2632 9367 2635
rect 10410 2632 10416 2644
rect 9355 2604 10416 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 12066 2632 12072 2644
rect 11931 2604 12072 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 15657 2635 15715 2641
rect 15657 2632 15669 2635
rect 12860 2604 15669 2632
rect 12860 2592 12866 2604
rect 15657 2601 15669 2604
rect 15703 2601 15715 2635
rect 15657 2595 15715 2601
rect 16206 2592 16212 2644
rect 16264 2592 16270 2644
rect 17034 2592 17040 2644
rect 17092 2592 17098 2644
rect 19518 2632 19524 2644
rect 17604 2604 19524 2632
rect 4982 2524 4988 2576
rect 5040 2524 5046 2576
rect 17604 2564 17632 2604
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 22833 2635 22891 2641
rect 22833 2601 22845 2635
rect 22879 2632 22891 2635
rect 23106 2632 23112 2644
rect 22879 2604 23112 2632
rect 22879 2601 22891 2604
rect 22833 2595 22891 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23290 2592 23296 2644
rect 23348 2632 23354 2644
rect 23385 2635 23443 2641
rect 23385 2632 23397 2635
rect 23348 2604 23397 2632
rect 23348 2592 23354 2604
rect 23385 2601 23397 2604
rect 23431 2601 23443 2635
rect 23385 2595 23443 2601
rect 23566 2592 23572 2644
rect 23624 2592 23630 2644
rect 23658 2592 23664 2644
rect 23716 2592 23722 2644
rect 6886 2536 17632 2564
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 5905 2499 5963 2505
rect 5905 2465 5917 2499
rect 5951 2496 5963 2499
rect 6886 2496 6914 2536
rect 17678 2524 17684 2576
rect 17736 2564 17742 2576
rect 20073 2567 20131 2573
rect 20073 2564 20085 2567
rect 17736 2536 20085 2564
rect 17736 2524 17742 2536
rect 20073 2533 20085 2536
rect 20119 2533 20131 2567
rect 20073 2527 20131 2533
rect 21174 2524 21180 2576
rect 21232 2564 21238 2576
rect 21232 2536 24900 2564
rect 21232 2524 21238 2536
rect 5951 2468 6914 2496
rect 7469 2499 7527 2505
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7515 2468 8248 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 992 2400 1777 2428
rect 992 2388 998 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 2004 2400 2053 2428
rect 2004 2388 2010 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4111 2400 5488 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4801 2363 4859 2369
rect 4801 2360 4813 2363
rect 4580 2332 4813 2360
rect 4580 2320 4586 2332
rect 4801 2329 4813 2332
rect 4847 2329 4859 2363
rect 5460 2360 5488 2400
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5868 2400 6193 2428
rect 5868 2388 5874 2400
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8113 2431 8171 2437
rect 7800 2424 8064 2428
rect 8113 2424 8125 2431
rect 7800 2400 8125 2424
rect 7800 2388 7806 2400
rect 8036 2397 8125 2400
rect 8159 2397 8171 2431
rect 8220 2428 8248 2468
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 10134 2496 10140 2508
rect 8352 2468 10140 2496
rect 8352 2456 8358 2468
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 10652 2468 11836 2496
rect 10652 2456 10658 2468
rect 8846 2428 8852 2440
rect 8220 2400 8852 2428
rect 8036 2396 8171 2397
rect 8113 2391 8171 2396
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10376 2400 10425 2428
rect 10376 2388 10382 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 11808 2428 11836 2468
rect 11882 2456 11888 2508
rect 11940 2496 11946 2508
rect 23658 2496 23664 2508
rect 11940 2468 23664 2496
rect 11940 2456 11946 2468
rect 23658 2456 23664 2468
rect 23716 2456 23722 2508
rect 24872 2505 24900 2536
rect 24857 2499 24915 2505
rect 24857 2465 24869 2499
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 12802 2428 12808 2440
rect 11808 2400 12808 2428
rect 10689 2391 10747 2397
rect 8938 2360 8944 2372
rect 5460 2332 8944 2360
rect 4801 2323 4859 2329
rect 8938 2320 8944 2332
rect 8996 2320 9002 2372
rect 1578 2252 1584 2304
rect 1636 2252 1642 2304
rect 1949 2295 2007 2301
rect 1949 2261 1961 2295
rect 1995 2292 2007 2295
rect 8018 2292 8024 2304
rect 1995 2264 8024 2292
rect 1995 2261 2007 2264
rect 1949 2255 2007 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 10704 2292 10732 2391
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12952 2400 13001 2428
rect 12952 2388 12958 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2428 14611 2431
rect 14599 2400 15884 2428
rect 14599 2397 14611 2400
rect 14553 2391 14611 2397
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 14182 2320 14188 2372
rect 14240 2360 14246 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 14240 2332 14381 2360
rect 14240 2320 14246 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 15470 2320 15476 2372
rect 15528 2360 15534 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 15528 2332 15761 2360
rect 15528 2320 15534 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 15856 2360 15884 2400
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16393 2431 16451 2437
rect 16393 2428 16405 2431
rect 16172 2400 16405 2428
rect 16172 2388 16178 2400
rect 16393 2397 16405 2400
rect 16439 2397 16451 2431
rect 16393 2391 16451 2397
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16540 2400 16957 2428
rect 16540 2388 16546 2400
rect 16945 2397 16957 2400
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 16574 2360 16580 2372
rect 15856 2332 16580 2360
rect 15749 2323 15807 2329
rect 16574 2320 16580 2332
rect 16632 2320 16638 2372
rect 16960 2360 16988 2391
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17460 2400 17509 2428
rect 17460 2388 17466 2400
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 19426 2428 19432 2440
rect 17497 2391 17555 2397
rect 17604 2400 19432 2428
rect 17604 2360 17632 2400
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 22554 2388 22560 2440
rect 22612 2428 22618 2440
rect 22649 2431 22707 2437
rect 22649 2428 22661 2431
rect 22612 2400 22661 2428
rect 22612 2388 22618 2400
rect 22649 2397 22661 2400
rect 22695 2397 22707 2431
rect 22649 2391 22707 2397
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23348 2400 23857 2428
rect 23348 2388 23354 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25866 2388 25872 2440
rect 25924 2388 25930 2440
rect 28445 2431 28503 2437
rect 28445 2428 28457 2431
rect 26206 2400 28457 2428
rect 16960 2332 17632 2360
rect 18690 2320 18696 2372
rect 18748 2360 18754 2372
rect 18969 2363 19027 2369
rect 18969 2360 18981 2363
rect 18748 2332 18981 2360
rect 18748 2320 18754 2332
rect 18969 2329 18981 2332
rect 19015 2329 19027 2363
rect 18969 2323 19027 2329
rect 19334 2320 19340 2372
rect 19392 2320 19398 2372
rect 23106 2320 23112 2372
rect 23164 2360 23170 2372
rect 23201 2363 23259 2369
rect 23201 2360 23213 2363
rect 23164 2332 23213 2360
rect 23164 2320 23170 2332
rect 23201 2329 23213 2332
rect 23247 2329 23259 2363
rect 23201 2323 23259 2329
rect 23382 2320 23388 2372
rect 23440 2369 23446 2372
rect 23440 2363 23459 2369
rect 23447 2329 23459 2363
rect 23440 2323 23459 2329
rect 23440 2320 23446 2323
rect 25774 2320 25780 2372
rect 25832 2360 25838 2372
rect 26053 2363 26111 2369
rect 26053 2360 26065 2363
rect 25832 2332 26065 2360
rect 25832 2320 25838 2332
rect 26053 2329 26065 2332
rect 26099 2329 26111 2363
rect 26053 2323 26111 2329
rect 15562 2292 15568 2304
rect 10704 2264 15568 2292
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 15654 2252 15660 2304
rect 15712 2292 15718 2304
rect 17727 2295 17785 2301
rect 17727 2292 17739 2295
rect 15712 2264 17739 2292
rect 15712 2252 15718 2264
rect 17727 2261 17739 2264
rect 17773 2261 17785 2295
rect 17727 2255 17785 2261
rect 18874 2252 18880 2304
rect 18932 2252 18938 2304
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 26206 2292 26234 2400
rect 28445 2397 28457 2400
rect 28491 2397 28503 2431
rect 29638 2428 29644 2440
rect 28445 2391 28503 2397
rect 29104 2400 29644 2428
rect 27062 2320 27068 2372
rect 27120 2360 27126 2372
rect 27341 2363 27399 2369
rect 27341 2360 27353 2363
rect 27120 2332 27353 2360
rect 27120 2320 27126 2332
rect 27341 2329 27353 2332
rect 27387 2329 27399 2363
rect 27341 2323 27399 2329
rect 28261 2363 28319 2369
rect 28261 2329 28273 2363
rect 28307 2329 28319 2363
rect 28261 2323 28319 2329
rect 20864 2264 26234 2292
rect 20864 2252 20870 2264
rect 27246 2252 27252 2304
rect 27304 2252 27310 2304
rect 28166 2252 28172 2304
rect 28224 2252 28230 2304
rect 28276 2292 28304 2323
rect 28350 2320 28356 2372
rect 28408 2360 28414 2372
rect 28629 2363 28687 2369
rect 28629 2360 28641 2363
rect 28408 2332 28641 2360
rect 28408 2320 28414 2332
rect 28629 2329 28641 2332
rect 28675 2329 28687 2363
rect 28629 2323 28687 2329
rect 29104 2292 29132 2400
rect 29638 2388 29644 2400
rect 29696 2388 29702 2440
rect 29270 2320 29276 2372
rect 29328 2320 29334 2372
rect 28276 2264 29132 2292
rect 29178 2252 29184 2304
rect 29236 2252 29242 2304
rect 1104 2202 29716 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 29716 2202
rect 1104 2128 29716 2150
rect 13998 1980 14004 2032
rect 14056 2020 14062 2032
rect 28166 2020 28172 2032
rect 14056 1992 28172 2020
rect 14056 1980 14062 1992
rect 28166 1980 28172 1992
rect 28224 1980 28230 2032
rect 1578 1912 1584 1964
rect 1636 1952 1642 1964
rect 21910 1952 21916 1964
rect 1636 1924 21916 1952
rect 1636 1912 1642 1924
rect 21910 1912 21916 1924
rect 21968 1912 21974 1964
rect 13262 1844 13268 1896
rect 13320 1884 13326 1896
rect 19610 1884 19616 1896
rect 13320 1856 19616 1884
rect 13320 1844 13326 1856
rect 19610 1844 19616 1856
rect 19668 1844 19674 1896
rect 11422 1776 11428 1828
rect 11480 1816 11486 1828
rect 27246 1816 27252 1828
rect 11480 1788 27252 1816
rect 11480 1776 11486 1788
rect 27246 1776 27252 1788
rect 27304 1776 27310 1828
rect 14458 1640 14464 1692
rect 14516 1680 14522 1692
rect 29178 1680 29184 1692
rect 14516 1652 29184 1680
rect 14516 1640 14522 1652
rect 29178 1640 29184 1652
rect 29236 1640 29242 1692
<< via1 >>
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 1308 30268 1360 30320
rect 2596 30268 2648 30320
rect 8392 30268 8444 30320
rect 9680 30268 9732 30320
rect 15476 30268 15528 30320
rect 19340 30268 19392 30320
rect 20628 30268 20680 30320
rect 21916 30268 21968 30320
rect 25136 30268 25188 30320
rect 27712 30268 27764 30320
rect 20 30200 72 30252
rect 848 30132 900 30184
rect 1952 30132 2004 30184
rect 3884 30200 3936 30252
rect 5264 30243 5316 30252
rect 5264 30209 5273 30243
rect 5273 30209 5307 30243
rect 5307 30209 5316 30243
rect 5264 30200 5316 30209
rect 7104 30200 7156 30252
rect 10968 30200 11020 30252
rect 12256 30200 12308 30252
rect 13544 30200 13596 30252
rect 14832 30200 14884 30252
rect 16764 30200 16816 30252
rect 18052 30200 18104 30252
rect 22560 30200 22612 30252
rect 23848 30200 23900 30252
rect 26424 30200 26476 30252
rect 30288 30268 30340 30320
rect 29368 30243 29420 30252
rect 29368 30209 29377 30243
rect 29377 30209 29411 30243
rect 29411 30209 29420 30243
rect 29368 30200 29420 30209
rect 2688 30064 2740 30116
rect 2964 30107 3016 30116
rect 2964 30073 2973 30107
rect 2973 30073 3007 30107
rect 3007 30073 3016 30107
rect 2964 30064 3016 30073
rect 3332 30107 3384 30116
rect 3332 30073 3341 30107
rect 3341 30073 3375 30107
rect 3375 30073 3384 30107
rect 3332 30064 3384 30073
rect 11612 30132 11664 30184
rect 16580 30132 16632 30184
rect 26516 30132 26568 30184
rect 29736 30132 29788 30184
rect 9496 30064 9548 30116
rect 12072 30064 12124 30116
rect 20720 30107 20772 30116
rect 20720 30073 20729 30107
rect 20729 30073 20763 30107
rect 20763 30073 20772 30107
rect 20720 30064 20772 30073
rect 22376 30064 22428 30116
rect 27804 30064 27856 30116
rect 5264 29996 5316 30048
rect 5448 30039 5500 30048
rect 5448 30005 5457 30039
rect 5457 30005 5491 30039
rect 5491 30005 5500 30039
rect 5448 29996 5500 30005
rect 12164 29996 12216 30048
rect 12532 30039 12584 30048
rect 12532 30005 12541 30039
rect 12541 30005 12575 30039
rect 12575 30005 12584 30039
rect 12532 29996 12584 30005
rect 13544 29996 13596 30048
rect 14924 29996 14976 30048
rect 15660 30039 15712 30048
rect 15660 30005 15669 30039
rect 15669 30005 15703 30039
rect 15703 30005 15712 30039
rect 15660 29996 15712 30005
rect 18328 30039 18380 30048
rect 18328 30005 18337 30039
rect 18337 30005 18371 30039
rect 18371 30005 18380 30039
rect 18328 29996 18380 30005
rect 19524 30039 19576 30048
rect 19524 30005 19533 30039
rect 19533 30005 19567 30039
rect 19567 30005 19576 30039
rect 19524 29996 19576 30005
rect 23940 29996 23992 30048
rect 24124 30039 24176 30048
rect 24124 30005 24133 30039
rect 24133 30005 24167 30039
rect 24167 30005 24176 30039
rect 24124 29996 24176 30005
rect 26148 29996 26200 30048
rect 28080 29996 28132 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 940 29656 992 29708
rect 9220 29588 9272 29640
rect 13544 29631 13596 29640
rect 13544 29597 13553 29631
rect 13553 29597 13587 29631
rect 13587 29597 13596 29631
rect 13544 29588 13596 29597
rect 28540 29631 28592 29640
rect 28540 29597 28549 29631
rect 28549 29597 28583 29631
rect 28583 29597 28592 29631
rect 28540 29588 28592 29597
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 29000 29588 29052 29640
rect 1216 29520 1268 29572
rect 2596 29563 2648 29572
rect 2596 29529 2605 29563
rect 2605 29529 2639 29563
rect 2639 29529 2648 29563
rect 2596 29520 2648 29529
rect 28356 29563 28408 29572
rect 28356 29529 28365 29563
rect 28365 29529 28399 29563
rect 28399 29529 28408 29563
rect 28356 29520 28408 29529
rect 28632 29520 28684 29572
rect 13084 29452 13136 29504
rect 29460 29452 29512 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 17868 29248 17920 29300
rect 15752 29180 15804 29232
rect 18788 29180 18840 29232
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 12440 29112 12492 29164
rect 13636 29112 13688 29164
rect 21088 29112 21140 29164
rect 29276 29155 29328 29164
rect 29276 29121 29285 29155
rect 29285 29121 29319 29155
rect 29319 29121 29328 29155
rect 29276 29112 29328 29121
rect 4712 29044 4764 29096
rect 12624 29044 12676 29096
rect 15476 29044 15528 29096
rect 11152 28976 11204 29028
rect 18052 29087 18104 29096
rect 18052 29053 18061 29087
rect 18061 29053 18095 29087
rect 18095 29053 18104 29087
rect 18052 29044 18104 29053
rect 14556 28908 14608 28960
rect 23480 28976 23532 29028
rect 29184 28976 29236 29028
rect 18512 28908 18564 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 5264 28704 5316 28756
rect 9312 28704 9364 28756
rect 15752 28704 15804 28756
rect 18788 28704 18840 28756
rect 7288 28543 7340 28552
rect 7288 28509 7297 28543
rect 7297 28509 7331 28543
rect 7331 28509 7340 28543
rect 7288 28500 7340 28509
rect 25320 28636 25372 28688
rect 10416 28568 10468 28620
rect 7564 28543 7616 28552
rect 7564 28509 7573 28543
rect 7573 28509 7607 28543
rect 7607 28509 7616 28543
rect 7564 28500 7616 28509
rect 7472 28364 7524 28416
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 12348 28500 12400 28552
rect 8024 28364 8076 28416
rect 9036 28407 9088 28416
rect 9036 28373 9045 28407
rect 9045 28373 9079 28407
rect 9079 28373 9088 28407
rect 9036 28364 9088 28373
rect 10508 28432 10560 28484
rect 11152 28432 11204 28484
rect 12716 28543 12768 28552
rect 12716 28509 12725 28543
rect 12725 28509 12759 28543
rect 12759 28509 12768 28543
rect 12716 28500 12768 28509
rect 13176 28500 13228 28552
rect 13636 28543 13688 28552
rect 13636 28509 13645 28543
rect 13645 28509 13679 28543
rect 13679 28509 13688 28543
rect 13636 28500 13688 28509
rect 16948 28500 17000 28552
rect 17408 28543 17460 28552
rect 17408 28509 17417 28543
rect 17417 28509 17451 28543
rect 17451 28509 17460 28543
rect 17408 28500 17460 28509
rect 18512 28568 18564 28620
rect 19984 28611 20036 28620
rect 19984 28577 19993 28611
rect 19993 28577 20027 28611
rect 20027 28577 20036 28611
rect 19984 28568 20036 28577
rect 17868 28543 17920 28552
rect 17868 28509 17885 28543
rect 17885 28509 17919 28543
rect 17919 28509 17920 28543
rect 17868 28500 17920 28509
rect 18236 28500 18288 28552
rect 14004 28432 14056 28484
rect 24032 28543 24084 28552
rect 24032 28509 24041 28543
rect 24041 28509 24075 28543
rect 24075 28509 24084 28543
rect 24032 28500 24084 28509
rect 24492 28500 24544 28552
rect 25504 28543 25556 28552
rect 25504 28509 25513 28543
rect 25513 28509 25547 28543
rect 25547 28509 25556 28543
rect 25504 28500 25556 28509
rect 27068 28543 27120 28552
rect 27068 28509 27077 28543
rect 27077 28509 27111 28543
rect 27111 28509 27120 28543
rect 27068 28500 27120 28509
rect 29092 28543 29144 28552
rect 29092 28509 29101 28543
rect 29101 28509 29135 28543
rect 29135 28509 29144 28543
rect 29092 28500 29144 28509
rect 11336 28364 11388 28416
rect 12900 28364 12952 28416
rect 13636 28364 13688 28416
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 17960 28364 18012 28416
rect 20260 28475 20312 28484
rect 20260 28441 20269 28475
rect 20269 28441 20303 28475
rect 20303 28441 20312 28475
rect 20260 28432 20312 28441
rect 21272 28432 21324 28484
rect 22008 28475 22060 28484
rect 22008 28441 22017 28475
rect 22017 28441 22051 28475
rect 22051 28441 22060 28475
rect 22008 28432 22060 28441
rect 23480 28432 23532 28484
rect 25780 28475 25832 28484
rect 25780 28441 25789 28475
rect 25789 28441 25823 28475
rect 25823 28441 25832 28475
rect 25780 28432 25832 28441
rect 27344 28475 27396 28484
rect 27344 28441 27353 28475
rect 27353 28441 27387 28475
rect 27387 28441 27396 28475
rect 27344 28432 27396 28441
rect 21088 28364 21140 28416
rect 24216 28364 24268 28416
rect 25964 28364 26016 28416
rect 27160 28364 27212 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 7288 28160 7340 28212
rect 4712 28024 4764 28076
rect 5908 28024 5960 28076
rect 6552 28067 6604 28076
rect 6552 28033 6561 28067
rect 6561 28033 6595 28067
rect 6595 28033 6604 28067
rect 6552 28024 6604 28033
rect 7104 27956 7156 28008
rect 5816 27820 5868 27872
rect 6460 27863 6512 27872
rect 6460 27829 6469 27863
rect 6469 27829 6503 27863
rect 6503 27829 6512 27863
rect 6460 27820 6512 27829
rect 8024 28135 8076 28144
rect 8024 28101 8033 28135
rect 8033 28101 8067 28135
rect 8067 28101 8076 28135
rect 8024 28092 8076 28101
rect 9036 28092 9088 28144
rect 10508 28203 10560 28212
rect 10508 28169 10517 28203
rect 10517 28169 10551 28203
rect 10551 28169 10560 28203
rect 10508 28160 10560 28169
rect 10692 28160 10744 28212
rect 12716 28160 12768 28212
rect 13176 28160 13228 28212
rect 13912 28160 13964 28212
rect 14556 28203 14608 28212
rect 14556 28169 14565 28203
rect 14565 28169 14599 28203
rect 14599 28169 14608 28203
rect 14556 28160 14608 28169
rect 14832 28160 14884 28212
rect 7748 27999 7800 28008
rect 7748 27965 7757 27999
rect 7757 27965 7791 27999
rect 7791 27965 7800 27999
rect 7748 27956 7800 27965
rect 7472 27888 7524 27940
rect 10048 28067 10100 28076
rect 10048 28033 10057 28067
rect 10057 28033 10091 28067
rect 10091 28033 10100 28067
rect 10048 28024 10100 28033
rect 10140 28067 10192 28076
rect 10140 28033 10149 28067
rect 10149 28033 10183 28067
rect 10183 28033 10192 28067
rect 10140 28024 10192 28033
rect 10232 28067 10284 28076
rect 10232 28033 10241 28067
rect 10241 28033 10275 28067
rect 10275 28033 10284 28067
rect 10232 28024 10284 28033
rect 12900 28135 12952 28144
rect 12900 28101 12909 28135
rect 12909 28101 12943 28135
rect 12943 28101 12952 28135
rect 12900 28092 12952 28101
rect 13636 28092 13688 28144
rect 14740 28135 14792 28144
rect 14740 28101 14749 28135
rect 14749 28101 14783 28135
rect 14783 28101 14792 28135
rect 14740 28092 14792 28101
rect 15292 28135 15344 28144
rect 15292 28101 15301 28135
rect 15301 28101 15335 28135
rect 15335 28101 15344 28135
rect 15292 28092 15344 28101
rect 11152 28067 11204 28076
rect 11152 28033 11161 28067
rect 11161 28033 11195 28067
rect 11195 28033 11204 28067
rect 11152 28024 11204 28033
rect 11336 28024 11388 28076
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 17408 28160 17460 28212
rect 17592 28160 17644 28212
rect 16120 28135 16172 28144
rect 16120 28101 16129 28135
rect 16129 28101 16163 28135
rect 16163 28101 16172 28135
rect 16120 28092 16172 28101
rect 19248 28160 19300 28212
rect 20260 28160 20312 28212
rect 21272 28160 21324 28212
rect 24492 28203 24544 28212
rect 24492 28169 24501 28203
rect 24501 28169 24535 28203
rect 24535 28169 24544 28203
rect 24492 28160 24544 28169
rect 17132 28024 17184 28076
rect 18512 28067 18564 28076
rect 18512 28033 18521 28067
rect 18521 28033 18555 28067
rect 18555 28033 18564 28067
rect 18512 28024 18564 28033
rect 19432 28092 19484 28144
rect 18972 28024 19024 28076
rect 22008 28092 22060 28144
rect 11060 27888 11112 27940
rect 12348 27888 12400 27940
rect 14188 27888 14240 27940
rect 15016 27888 15068 27940
rect 21088 27956 21140 28008
rect 23480 28067 23532 28076
rect 23480 28033 23489 28067
rect 23489 28033 23523 28067
rect 23523 28033 23532 28067
rect 23480 28024 23532 28033
rect 24216 28067 24268 28076
rect 24216 28033 24225 28067
rect 24225 28033 24259 28067
rect 24259 28033 24268 28067
rect 25136 28092 25188 28144
rect 29092 28092 29144 28144
rect 24216 28024 24268 28033
rect 27160 28067 27212 28076
rect 27160 28033 27169 28067
rect 27169 28033 27203 28067
rect 27203 28033 27212 28067
rect 27160 28024 27212 28033
rect 23664 27956 23716 28008
rect 24032 27956 24084 28008
rect 24768 27999 24820 28008
rect 24768 27965 24777 27999
rect 24777 27965 24811 27999
rect 24811 27965 24820 27999
rect 24768 27956 24820 27965
rect 25044 27999 25096 28008
rect 25044 27965 25053 27999
rect 25053 27965 25087 27999
rect 25087 27965 25096 27999
rect 25044 27956 25096 27965
rect 25780 27956 25832 28008
rect 9128 27820 9180 27872
rect 10784 27863 10836 27872
rect 10784 27829 10793 27863
rect 10793 27829 10827 27863
rect 10827 27829 10836 27863
rect 10784 27820 10836 27829
rect 14648 27820 14700 27872
rect 15476 27863 15528 27872
rect 15476 27829 15485 27863
rect 15485 27829 15519 27863
rect 15519 27829 15528 27863
rect 15476 27820 15528 27829
rect 16396 27820 16448 27872
rect 16764 27863 16816 27872
rect 16764 27829 16773 27863
rect 16773 27829 16807 27863
rect 16807 27829 16816 27863
rect 16764 27820 16816 27829
rect 17868 27820 17920 27872
rect 19432 27820 19484 27872
rect 23848 27863 23900 27872
rect 23848 27829 23857 27863
rect 23857 27829 23891 27863
rect 23891 27829 23900 27863
rect 23848 27820 23900 27829
rect 25504 27820 25556 27872
rect 27344 27956 27396 28008
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 10048 27616 10100 27668
rect 10784 27616 10836 27668
rect 14188 27659 14240 27668
rect 14188 27625 14197 27659
rect 14197 27625 14231 27659
rect 14231 27625 14240 27659
rect 14188 27616 14240 27625
rect 14740 27616 14792 27668
rect 16120 27616 16172 27668
rect 16396 27616 16448 27668
rect 17868 27659 17920 27668
rect 17868 27625 17877 27659
rect 17877 27625 17911 27659
rect 17911 27625 17920 27659
rect 17868 27616 17920 27625
rect 18052 27659 18104 27668
rect 18052 27625 18061 27659
rect 18061 27625 18095 27659
rect 18095 27625 18104 27659
rect 18052 27616 18104 27625
rect 6368 27548 6420 27600
rect 6552 27591 6604 27600
rect 6552 27557 6561 27591
rect 6561 27557 6595 27591
rect 6595 27557 6604 27591
rect 6552 27548 6604 27557
rect 3700 27480 3752 27532
rect 4804 27523 4856 27532
rect 4804 27489 4813 27523
rect 4813 27489 4847 27523
rect 4847 27489 4856 27523
rect 4804 27480 4856 27489
rect 848 27412 900 27464
rect 1676 27455 1728 27464
rect 1676 27421 1685 27455
rect 1685 27421 1719 27455
rect 1719 27421 1728 27455
rect 1676 27412 1728 27421
rect 6460 27412 6512 27464
rect 6828 27412 6880 27464
rect 7380 27455 7432 27464
rect 7380 27421 7389 27455
rect 7389 27421 7423 27455
rect 7423 27421 7432 27455
rect 7380 27412 7432 27421
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 10692 27591 10744 27600
rect 10692 27557 10701 27591
rect 10701 27557 10735 27591
rect 10735 27557 10744 27591
rect 10692 27548 10744 27557
rect 13176 27591 13228 27600
rect 13176 27557 13185 27591
rect 13185 27557 13219 27591
rect 13219 27557 13228 27591
rect 13176 27548 13228 27557
rect 17132 27548 17184 27600
rect 17592 27548 17644 27600
rect 17776 27548 17828 27600
rect 18972 27616 19024 27668
rect 19432 27616 19484 27668
rect 23848 27616 23900 27668
rect 25044 27616 25096 27668
rect 25780 27659 25832 27668
rect 25780 27625 25789 27659
rect 25789 27625 25823 27659
rect 25823 27625 25832 27659
rect 25780 27616 25832 27625
rect 19616 27548 19668 27600
rect 8208 27480 8260 27532
rect 8484 27412 8536 27464
rect 9128 27455 9180 27464
rect 9128 27421 9137 27455
rect 9137 27421 9171 27455
rect 9171 27421 9180 27455
rect 9128 27412 9180 27421
rect 10140 27480 10192 27532
rect 10048 27455 10100 27464
rect 10048 27421 10057 27455
rect 10057 27421 10091 27455
rect 10091 27421 10100 27455
rect 10048 27412 10100 27421
rect 10232 27412 10284 27464
rect 11336 27455 11388 27464
rect 11336 27421 11345 27455
rect 11345 27421 11379 27455
rect 11379 27421 11388 27455
rect 11336 27412 11388 27421
rect 15016 27480 15068 27532
rect 14004 27412 14056 27464
rect 14372 27455 14424 27464
rect 14372 27421 14381 27455
rect 14381 27421 14415 27455
rect 14415 27421 14424 27455
rect 14372 27412 14424 27421
rect 5356 27344 5408 27396
rect 5816 27344 5868 27396
rect 6368 27344 6420 27396
rect 7104 27387 7156 27396
rect 7104 27353 7113 27387
rect 7113 27353 7147 27387
rect 7147 27353 7156 27387
rect 7104 27344 7156 27353
rect 7840 27387 7892 27396
rect 7840 27353 7849 27387
rect 7849 27353 7883 27387
rect 7883 27353 7892 27387
rect 7840 27344 7892 27353
rect 8024 27344 8076 27396
rect 10968 27344 11020 27396
rect 11060 27387 11112 27396
rect 11060 27353 11069 27387
rect 11069 27353 11103 27387
rect 11103 27353 11112 27387
rect 11060 27344 11112 27353
rect 6644 27276 6696 27328
rect 7656 27319 7708 27328
rect 7656 27285 7665 27319
rect 7665 27285 7699 27319
rect 7699 27285 7708 27319
rect 7656 27276 7708 27285
rect 8116 27319 8168 27328
rect 8116 27285 8125 27319
rect 8125 27285 8159 27319
rect 8159 27285 8168 27319
rect 8116 27276 8168 27285
rect 9128 27276 9180 27328
rect 12624 27344 12676 27396
rect 14096 27344 14148 27396
rect 14832 27412 14884 27464
rect 15384 27412 15436 27464
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 19984 27480 20036 27532
rect 23480 27480 23532 27532
rect 15292 27344 15344 27396
rect 15568 27344 15620 27396
rect 16764 27344 16816 27396
rect 17960 27344 18012 27396
rect 19248 27455 19300 27464
rect 19248 27421 19257 27455
rect 19257 27421 19291 27455
rect 19291 27421 19300 27455
rect 19248 27412 19300 27421
rect 19708 27412 19760 27464
rect 24768 27412 24820 27464
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 25320 27455 25372 27464
rect 25320 27421 25329 27455
rect 25329 27421 25363 27455
rect 25363 27421 25372 27455
rect 25320 27412 25372 27421
rect 27068 27412 27120 27464
rect 27620 27455 27672 27464
rect 27620 27421 27629 27455
rect 27629 27421 27663 27455
rect 27663 27421 27672 27455
rect 27620 27412 27672 27421
rect 13268 27276 13320 27328
rect 13544 27276 13596 27328
rect 14188 27276 14240 27328
rect 14372 27276 14424 27328
rect 19340 27276 19392 27328
rect 21180 27344 21232 27396
rect 22560 27344 22612 27396
rect 20628 27276 20680 27328
rect 25504 27344 25556 27396
rect 25872 27344 25924 27396
rect 25964 27387 26016 27396
rect 25964 27353 25973 27387
rect 25973 27353 26007 27387
rect 26007 27353 26016 27387
rect 25964 27344 26016 27353
rect 27896 27387 27948 27396
rect 27896 27353 27905 27387
rect 27905 27353 27939 27387
rect 27939 27353 27948 27387
rect 27896 27344 27948 27353
rect 28908 27344 28960 27396
rect 27988 27276 28040 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 5356 27072 5408 27124
rect 6644 27072 6696 27124
rect 7564 27072 7616 27124
rect 8484 27072 8536 27124
rect 9588 27115 9640 27124
rect 9588 27081 9597 27115
rect 9597 27081 9631 27115
rect 9631 27081 9640 27115
rect 9588 27072 9640 27081
rect 12624 27072 12676 27124
rect 14004 27115 14056 27124
rect 14004 27081 14013 27115
rect 14013 27081 14047 27115
rect 14047 27081 14056 27115
rect 14004 27072 14056 27081
rect 18512 27072 18564 27124
rect 19340 27072 19392 27124
rect 20628 27072 20680 27124
rect 21180 27072 21232 27124
rect 22560 27072 22612 27124
rect 27896 27072 27948 27124
rect 28908 27115 28960 27124
rect 28908 27081 28917 27115
rect 28917 27081 28951 27115
rect 28951 27081 28960 27115
rect 28908 27072 28960 27081
rect 6184 27004 6236 27056
rect 6828 27004 6880 27056
rect 6920 26979 6972 26988
rect 6920 26945 6929 26979
rect 6929 26945 6963 26979
rect 6963 26945 6972 26979
rect 6920 26936 6972 26945
rect 7288 27004 7340 27056
rect 8024 27004 8076 27056
rect 8116 27047 8168 27056
rect 8116 27013 8125 27047
rect 8125 27013 8159 27047
rect 8159 27013 8168 27047
rect 8116 27004 8168 27013
rect 9128 27004 9180 27056
rect 7748 26936 7800 26988
rect 7380 26868 7432 26920
rect 10324 26868 10376 26920
rect 3332 26800 3384 26852
rect 19248 27004 19300 27056
rect 24492 27004 24544 27056
rect 29276 27047 29328 27056
rect 29276 27013 29285 27047
rect 29285 27013 29319 27047
rect 29319 27013 29328 27047
rect 29276 27004 29328 27013
rect 10968 26936 11020 26988
rect 12440 26936 12492 26988
rect 13268 26979 13320 26988
rect 13268 26945 13277 26979
rect 13277 26945 13311 26979
rect 13311 26945 13320 26979
rect 13268 26936 13320 26945
rect 14096 26979 14148 26988
rect 14096 26945 14105 26979
rect 14105 26945 14139 26979
rect 14139 26945 14148 26979
rect 14096 26936 14148 26945
rect 14832 26979 14884 26988
rect 14832 26945 14841 26979
rect 14841 26945 14875 26979
rect 14875 26945 14884 26979
rect 14832 26936 14884 26945
rect 15936 26936 15988 26988
rect 18604 26936 18656 26988
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 21088 26936 21140 26988
rect 22008 26936 22060 26988
rect 11152 26868 11204 26920
rect 13728 26868 13780 26920
rect 23480 26868 23532 26920
rect 23756 26868 23808 26920
rect 24952 26911 25004 26920
rect 24952 26877 24961 26911
rect 24961 26877 24995 26911
rect 24995 26877 25004 26911
rect 24952 26868 25004 26877
rect 6828 26732 6880 26784
rect 6920 26732 6972 26784
rect 7380 26732 7432 26784
rect 12624 26800 12676 26852
rect 13452 26800 13504 26852
rect 17868 26800 17920 26852
rect 18420 26800 18472 26852
rect 20720 26800 20772 26852
rect 10048 26732 10100 26784
rect 13176 26732 13228 26784
rect 13544 26732 13596 26784
rect 15200 26775 15252 26784
rect 15200 26741 15209 26775
rect 15209 26741 15243 26775
rect 15243 26741 15252 26775
rect 15200 26732 15252 26741
rect 15292 26732 15344 26784
rect 15752 26732 15804 26784
rect 23480 26775 23532 26784
rect 23480 26741 23489 26775
rect 23489 26741 23523 26775
rect 23523 26741 23532 26775
rect 23480 26732 23532 26741
rect 24768 26732 24820 26784
rect 27068 26936 27120 26988
rect 27988 26936 28040 26988
rect 29092 26936 29144 26988
rect 27436 26911 27488 26920
rect 27436 26877 27445 26911
rect 27445 26877 27479 26911
rect 27479 26877 27488 26911
rect 27436 26868 27488 26877
rect 29552 26732 29604 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 4804 26392 4856 26444
rect 4712 26367 4764 26376
rect 1492 26299 1544 26308
rect 1492 26265 1501 26299
rect 1501 26265 1535 26299
rect 1535 26265 1544 26299
rect 1492 26256 1544 26265
rect 2044 26256 2096 26308
rect 4160 26256 4212 26308
rect 4712 26333 4721 26367
rect 4721 26333 4755 26367
rect 4755 26333 4764 26367
rect 4712 26324 4764 26333
rect 16856 26528 16908 26580
rect 12624 26460 12676 26512
rect 8484 26392 8536 26444
rect 4620 26231 4672 26240
rect 4620 26197 4629 26231
rect 4629 26197 4663 26231
rect 4663 26197 4672 26231
rect 4620 26188 4672 26197
rect 4712 26188 4764 26240
rect 5264 26256 5316 26308
rect 6000 26299 6052 26308
rect 6000 26265 6009 26299
rect 6009 26265 6043 26299
rect 6043 26265 6052 26299
rect 6000 26256 6052 26265
rect 6644 26324 6696 26376
rect 8576 26324 8628 26376
rect 9404 26367 9456 26376
rect 9404 26333 9413 26367
rect 9413 26333 9447 26367
rect 9447 26333 9456 26367
rect 9404 26324 9456 26333
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 10324 26367 10376 26376
rect 10324 26333 10333 26367
rect 10333 26333 10367 26367
rect 10367 26333 10376 26367
rect 10324 26324 10376 26333
rect 11244 26324 11296 26376
rect 11704 26392 11756 26444
rect 13176 26435 13228 26444
rect 13176 26401 13185 26435
rect 13185 26401 13219 26435
rect 13219 26401 13228 26435
rect 13176 26392 13228 26401
rect 5356 26188 5408 26240
rect 6276 26188 6328 26240
rect 6460 26188 6512 26240
rect 6736 26188 6788 26240
rect 7196 26188 7248 26240
rect 7656 26188 7708 26240
rect 8300 26231 8352 26240
rect 8300 26197 8309 26231
rect 8309 26197 8343 26231
rect 8343 26197 8352 26231
rect 8300 26188 8352 26197
rect 9864 26188 9916 26240
rect 10600 26299 10652 26308
rect 10600 26265 10609 26299
rect 10609 26265 10643 26299
rect 10643 26265 10652 26299
rect 10600 26256 10652 26265
rect 10876 26256 10928 26308
rect 12900 26367 12952 26376
rect 12900 26333 12909 26367
rect 12909 26333 12943 26367
rect 12943 26333 12952 26367
rect 12900 26324 12952 26333
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 13084 26367 13136 26376
rect 13084 26333 13093 26367
rect 13093 26333 13127 26367
rect 13127 26333 13136 26367
rect 13084 26324 13136 26333
rect 14648 26435 14700 26444
rect 14648 26401 14657 26435
rect 14657 26401 14691 26435
rect 14691 26401 14700 26435
rect 14648 26392 14700 26401
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 15752 26324 15804 26376
rect 17132 26460 17184 26512
rect 23296 26460 23348 26512
rect 23756 26571 23808 26580
rect 23756 26537 23765 26571
rect 23765 26537 23799 26571
rect 23799 26537 23808 26571
rect 23756 26528 23808 26537
rect 24952 26528 25004 26580
rect 17224 26435 17276 26444
rect 17224 26401 17233 26435
rect 17233 26401 17267 26435
rect 17267 26401 17276 26435
rect 17224 26392 17276 26401
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 10968 26231 11020 26240
rect 10968 26197 10977 26231
rect 10977 26197 11011 26231
rect 11011 26197 11020 26231
rect 10968 26188 11020 26197
rect 12440 26231 12492 26240
rect 12440 26197 12449 26231
rect 12449 26197 12483 26231
rect 12483 26197 12492 26231
rect 12440 26188 12492 26197
rect 12716 26188 12768 26240
rect 13636 26231 13688 26240
rect 13636 26197 13645 26231
rect 13645 26197 13679 26231
rect 13679 26197 13688 26231
rect 13636 26188 13688 26197
rect 16212 26299 16264 26308
rect 16212 26265 16221 26299
rect 16221 26265 16255 26299
rect 16255 26265 16264 26299
rect 16212 26256 16264 26265
rect 18052 26324 18104 26376
rect 17684 26299 17736 26308
rect 17684 26265 17693 26299
rect 17693 26265 17727 26299
rect 17727 26265 17736 26299
rect 17684 26256 17736 26265
rect 18144 26256 18196 26308
rect 18420 26324 18472 26376
rect 18604 26367 18656 26376
rect 18604 26333 18613 26367
rect 18613 26333 18647 26367
rect 18647 26333 18656 26367
rect 18604 26324 18656 26333
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 18972 26367 19024 26376
rect 18972 26333 18981 26367
rect 18981 26333 19015 26367
rect 19015 26333 19024 26367
rect 18972 26324 19024 26333
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 16396 26188 16448 26240
rect 18788 26299 18840 26308
rect 18788 26265 18797 26299
rect 18797 26265 18831 26299
rect 18831 26265 18840 26299
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 20076 26367 20128 26376
rect 20076 26333 20085 26367
rect 20085 26333 20119 26367
rect 20119 26333 20128 26367
rect 20076 26324 20128 26333
rect 18788 26256 18840 26265
rect 20260 26256 20312 26308
rect 19340 26188 19392 26240
rect 19800 26231 19852 26240
rect 19800 26197 19809 26231
rect 19809 26197 19843 26231
rect 19843 26197 19852 26231
rect 19800 26188 19852 26197
rect 23388 26324 23440 26376
rect 24768 26392 24820 26444
rect 25872 26392 25924 26444
rect 27988 26503 28040 26512
rect 27988 26469 27997 26503
rect 27997 26469 28031 26503
rect 28031 26469 28040 26503
rect 27988 26460 28040 26469
rect 21824 26188 21876 26240
rect 23480 26299 23532 26308
rect 23480 26265 23489 26299
rect 23489 26265 23523 26299
rect 23523 26265 23532 26299
rect 23480 26256 23532 26265
rect 23664 26256 23716 26308
rect 26976 26367 27028 26376
rect 26976 26333 26985 26367
rect 26985 26333 27019 26367
rect 27019 26333 27028 26367
rect 26976 26324 27028 26333
rect 25228 26299 25280 26308
rect 25228 26265 25237 26299
rect 25237 26265 25271 26299
rect 25271 26265 25280 26299
rect 25228 26256 25280 26265
rect 26240 26256 26292 26308
rect 23940 26231 23992 26240
rect 23940 26197 23949 26231
rect 23949 26197 23983 26231
rect 23983 26197 23992 26231
rect 23940 26188 23992 26197
rect 26792 26231 26844 26240
rect 26792 26197 26801 26231
rect 26801 26197 26835 26231
rect 26835 26197 26844 26231
rect 26792 26188 26844 26197
rect 27344 26324 27396 26376
rect 29276 26299 29328 26308
rect 29276 26265 29285 26299
rect 29285 26265 29319 26299
rect 29319 26265 29328 26299
rect 29276 26256 29328 26265
rect 27344 26188 27396 26240
rect 27804 26231 27856 26240
rect 27804 26197 27813 26231
rect 27813 26197 27847 26231
rect 27847 26197 27856 26231
rect 27804 26188 27856 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 2596 25984 2648 26036
rect 5356 25984 5408 26036
rect 6000 25984 6052 26036
rect 6736 25984 6788 26036
rect 4712 25916 4764 25968
rect 6092 25916 6144 25968
rect 3700 25891 3752 25900
rect 3700 25857 3709 25891
rect 3709 25857 3743 25891
rect 3743 25857 3752 25891
rect 3700 25848 3752 25857
rect 5724 25848 5776 25900
rect 3976 25823 4028 25832
rect 3976 25789 3985 25823
rect 3985 25789 4019 25823
rect 4019 25789 4028 25823
rect 3976 25780 4028 25789
rect 6276 25848 6328 25900
rect 6644 25891 6696 25900
rect 6644 25857 6653 25891
rect 6653 25857 6687 25891
rect 6687 25857 6696 25891
rect 6644 25848 6696 25857
rect 8300 25916 8352 25968
rect 6920 25848 6972 25900
rect 7564 25891 7616 25900
rect 7564 25857 7573 25891
rect 7573 25857 7607 25891
rect 7607 25857 7616 25891
rect 7564 25848 7616 25857
rect 7748 25891 7800 25900
rect 7748 25857 7755 25891
rect 7755 25857 7800 25891
rect 7748 25848 7800 25857
rect 7840 25891 7892 25900
rect 7840 25857 7849 25891
rect 7849 25857 7883 25891
rect 7883 25857 7892 25891
rect 7840 25848 7892 25857
rect 6552 25712 6604 25764
rect 7472 25780 7524 25832
rect 7012 25712 7064 25764
rect 8392 25712 8444 25764
rect 7104 25644 7156 25696
rect 7656 25644 7708 25696
rect 7932 25644 7984 25696
rect 9220 25891 9272 25900
rect 9220 25857 9229 25891
rect 9229 25857 9263 25891
rect 9263 25857 9272 25891
rect 9220 25848 9272 25857
rect 10876 25984 10928 26036
rect 9864 25891 9916 25900
rect 9864 25857 9873 25891
rect 9873 25857 9907 25891
rect 9907 25857 9916 25891
rect 9864 25848 9916 25857
rect 9772 25780 9824 25832
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 10968 25891 11020 25900
rect 10968 25857 10977 25891
rect 10977 25857 11011 25891
rect 11011 25857 11020 25891
rect 12440 25984 12492 26036
rect 13636 25984 13688 26036
rect 14832 25984 14884 26036
rect 15200 26027 15252 26036
rect 15200 25993 15209 26027
rect 15209 25993 15243 26027
rect 15243 25993 15252 26027
rect 15200 25984 15252 25993
rect 10968 25848 11020 25857
rect 11888 25848 11940 25900
rect 12256 25891 12308 25900
rect 12256 25857 12265 25891
rect 12265 25857 12299 25891
rect 12299 25857 12308 25891
rect 12256 25848 12308 25857
rect 12900 25848 12952 25900
rect 9404 25712 9456 25764
rect 9864 25712 9916 25764
rect 9956 25687 10008 25696
rect 9956 25653 9965 25687
rect 9965 25653 9999 25687
rect 9999 25653 10008 25687
rect 9956 25644 10008 25653
rect 12624 25687 12676 25696
rect 12624 25653 12633 25687
rect 12633 25653 12667 25687
rect 12667 25653 12676 25687
rect 12624 25644 12676 25653
rect 12808 25712 12860 25764
rect 13084 25823 13136 25832
rect 13084 25789 13093 25823
rect 13093 25789 13127 25823
rect 13127 25789 13136 25823
rect 13084 25780 13136 25789
rect 13360 25891 13412 25900
rect 13360 25857 13369 25891
rect 13369 25857 13403 25891
rect 13403 25857 13412 25891
rect 13360 25848 13412 25857
rect 13452 25848 13504 25900
rect 13912 25848 13964 25900
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 15016 25916 15068 25968
rect 14280 25780 14332 25832
rect 14832 25823 14884 25832
rect 14832 25789 14841 25823
rect 14841 25789 14875 25823
rect 14875 25789 14884 25823
rect 14832 25780 14884 25789
rect 13176 25644 13228 25696
rect 13452 25644 13504 25696
rect 14464 25644 14516 25696
rect 14832 25644 14884 25696
rect 15752 25984 15804 26036
rect 15936 26027 15988 26036
rect 15936 25993 15945 26027
rect 15945 25993 15979 26027
rect 15979 25993 15988 26027
rect 15936 25984 15988 25993
rect 16212 25984 16264 26036
rect 18604 25984 18656 26036
rect 17040 25959 17092 25968
rect 17040 25925 17049 25959
rect 17049 25925 17083 25959
rect 17083 25925 17092 25959
rect 17040 25916 17092 25925
rect 17684 25916 17736 25968
rect 18972 25916 19024 25968
rect 15844 25848 15896 25900
rect 16212 25780 16264 25832
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17868 25848 17920 25900
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 18144 25891 18196 25900
rect 18144 25857 18153 25891
rect 18153 25857 18187 25891
rect 18187 25857 18196 25891
rect 18144 25848 18196 25857
rect 18420 25891 18472 25900
rect 18420 25857 18429 25891
rect 18429 25857 18463 25891
rect 18463 25857 18472 25891
rect 18420 25848 18472 25857
rect 21824 26027 21876 26036
rect 21824 25993 21833 26027
rect 21833 25993 21867 26027
rect 21867 25993 21876 26027
rect 21824 25984 21876 25993
rect 24492 25984 24544 26036
rect 25228 25984 25280 26036
rect 26240 25984 26292 26036
rect 27804 25984 27856 26036
rect 19432 25916 19484 25968
rect 20260 25916 20312 25968
rect 21456 25916 21508 25968
rect 22284 25916 22336 25968
rect 23296 25959 23348 25968
rect 23296 25925 23305 25959
rect 23305 25925 23339 25959
rect 23339 25925 23348 25959
rect 23296 25916 23348 25925
rect 25872 25916 25924 25968
rect 27344 25959 27396 25968
rect 27344 25925 27353 25959
rect 27353 25925 27387 25959
rect 27387 25925 27396 25959
rect 27344 25916 27396 25925
rect 17592 25780 17644 25832
rect 18788 25712 18840 25764
rect 16396 25687 16448 25696
rect 16396 25653 16405 25687
rect 16405 25653 16439 25687
rect 16439 25653 16448 25687
rect 16396 25644 16448 25653
rect 17408 25644 17460 25696
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 19892 25891 19944 25900
rect 19892 25857 19901 25891
rect 19901 25857 19935 25891
rect 19935 25857 19944 25891
rect 19892 25848 19944 25857
rect 24768 25848 24820 25900
rect 26240 25891 26292 25900
rect 22008 25780 22060 25832
rect 26240 25857 26249 25891
rect 26249 25857 26283 25891
rect 26283 25857 26292 25891
rect 26240 25848 26292 25857
rect 27160 25891 27212 25900
rect 27160 25857 27169 25891
rect 27169 25857 27203 25891
rect 27203 25857 27212 25891
rect 27160 25848 27212 25857
rect 29000 25848 29052 25900
rect 27620 25823 27672 25832
rect 27620 25789 27629 25823
rect 27629 25789 27663 25823
rect 27663 25789 27672 25823
rect 27620 25780 27672 25789
rect 27988 25780 28040 25832
rect 19432 25712 19484 25764
rect 26792 25712 26844 25764
rect 27712 25644 27764 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 3976 25440 4028 25492
rect 4620 25440 4672 25492
rect 9220 25440 9272 25492
rect 9680 25440 9732 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 11888 25483 11940 25492
rect 11888 25449 11897 25483
rect 11897 25449 11931 25483
rect 11931 25449 11940 25483
rect 11888 25440 11940 25449
rect 12992 25440 13044 25492
rect 13360 25440 13412 25492
rect 14464 25483 14516 25492
rect 14464 25449 14473 25483
rect 14473 25449 14507 25483
rect 14507 25449 14516 25483
rect 14464 25440 14516 25449
rect 16948 25440 17000 25492
rect 17592 25483 17644 25492
rect 17592 25449 17601 25483
rect 17601 25449 17635 25483
rect 17635 25449 17644 25483
rect 17592 25440 17644 25449
rect 18420 25440 18472 25492
rect 21456 25483 21508 25492
rect 21456 25449 21465 25483
rect 21465 25449 21499 25483
rect 21499 25449 21508 25483
rect 21456 25440 21508 25449
rect 22284 25483 22336 25492
rect 22284 25449 22293 25483
rect 22293 25449 22327 25483
rect 22327 25449 22336 25483
rect 22284 25440 22336 25449
rect 27436 25440 27488 25492
rect 27988 25483 28040 25492
rect 27988 25449 27997 25483
rect 27997 25449 28031 25483
rect 28031 25449 28040 25483
rect 27988 25440 28040 25449
rect 29000 25440 29052 25492
rect 6276 25372 6328 25424
rect 7932 25372 7984 25424
rect 10692 25372 10744 25424
rect 12256 25372 12308 25424
rect 13084 25372 13136 25424
rect 17040 25372 17092 25424
rect 4712 25279 4764 25288
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 5908 25236 5960 25288
rect 6000 25236 6052 25288
rect 6368 25279 6420 25288
rect 6368 25245 6375 25279
rect 6375 25245 6420 25279
rect 6368 25236 6420 25245
rect 6736 25236 6788 25288
rect 7196 25279 7248 25288
rect 7196 25245 7205 25279
rect 7205 25245 7239 25279
rect 7239 25245 7248 25279
rect 7196 25236 7248 25245
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 7656 25279 7708 25288
rect 7656 25245 7665 25279
rect 7665 25245 7699 25279
rect 7699 25245 7708 25279
rect 7656 25236 7708 25245
rect 6460 25211 6512 25220
rect 6460 25177 6469 25211
rect 6469 25177 6503 25211
rect 6503 25177 6512 25211
rect 6460 25168 6512 25177
rect 8024 25168 8076 25220
rect 8392 25304 8444 25356
rect 8668 25279 8720 25288
rect 8668 25245 8677 25279
rect 8677 25245 8711 25279
rect 8711 25245 8720 25279
rect 8668 25236 8720 25245
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9680 25236 9732 25245
rect 9772 25279 9824 25288
rect 9772 25245 9781 25279
rect 9781 25245 9815 25279
rect 9815 25245 9824 25279
rect 9772 25236 9824 25245
rect 10600 25236 10652 25288
rect 10692 25236 10744 25288
rect 10416 25168 10468 25220
rect 11244 25304 11296 25356
rect 11152 25279 11204 25288
rect 11152 25245 11161 25279
rect 11161 25245 11195 25279
rect 11195 25245 11204 25279
rect 11152 25236 11204 25245
rect 12900 25236 12952 25288
rect 13268 25304 13320 25356
rect 13452 25279 13504 25288
rect 13452 25245 13461 25279
rect 13461 25245 13495 25279
rect 13495 25245 13504 25279
rect 13452 25236 13504 25245
rect 17868 25304 17920 25356
rect 19708 25304 19760 25356
rect 20536 25304 20588 25356
rect 3884 25100 3936 25152
rect 6184 25100 6236 25152
rect 6828 25143 6880 25152
rect 6828 25109 6837 25143
rect 6837 25109 6871 25143
rect 6871 25109 6880 25143
rect 6828 25100 6880 25109
rect 7380 25143 7432 25152
rect 7380 25109 7389 25143
rect 7389 25109 7423 25143
rect 7423 25109 7432 25143
rect 7380 25100 7432 25109
rect 8116 25100 8168 25152
rect 9772 25100 9824 25152
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 13268 25211 13320 25220
rect 13268 25177 13277 25211
rect 13277 25177 13311 25211
rect 13311 25177 13320 25211
rect 13268 25168 13320 25177
rect 13636 25168 13688 25220
rect 12348 25100 12400 25152
rect 14280 25236 14332 25288
rect 15844 25279 15896 25288
rect 15844 25245 15853 25279
rect 15853 25245 15887 25279
rect 15887 25245 15896 25279
rect 15844 25236 15896 25245
rect 16672 25236 16724 25288
rect 17040 25279 17092 25288
rect 17040 25245 17049 25279
rect 17049 25245 17083 25279
rect 17083 25245 17092 25279
rect 17040 25236 17092 25245
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 18512 25236 18564 25288
rect 20076 25236 20128 25288
rect 22008 25236 22060 25288
rect 23572 25236 23624 25288
rect 23756 25236 23808 25288
rect 26792 25236 26844 25288
rect 27160 25236 27212 25288
rect 27344 25236 27396 25288
rect 27712 25236 27764 25288
rect 14188 25211 14240 25220
rect 14188 25177 14197 25211
rect 14197 25177 14231 25211
rect 14231 25177 14240 25211
rect 14188 25168 14240 25177
rect 26240 25168 26292 25220
rect 29092 25236 29144 25288
rect 14648 25100 14700 25152
rect 15936 25100 15988 25152
rect 19524 25100 19576 25152
rect 19800 25143 19852 25152
rect 19800 25109 19809 25143
rect 19809 25109 19843 25143
rect 19843 25109 19852 25143
rect 19800 25100 19852 25109
rect 23112 25100 23164 25152
rect 24032 25100 24084 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 5172 24896 5224 24948
rect 5356 24896 5408 24948
rect 5632 24939 5684 24948
rect 5632 24905 5641 24939
rect 5641 24905 5675 24939
rect 5675 24905 5684 24939
rect 5632 24896 5684 24905
rect 5908 24896 5960 24948
rect 6828 24896 6880 24948
rect 7104 24896 7156 24948
rect 14280 24896 14332 24948
rect 15844 24896 15896 24948
rect 16672 24939 16724 24948
rect 16672 24905 16681 24939
rect 16681 24905 16715 24939
rect 16715 24905 16724 24939
rect 16672 24896 16724 24905
rect 16856 24896 16908 24948
rect 848 24760 900 24812
rect 5356 24760 5408 24812
rect 5724 24760 5776 24812
rect 6644 24760 6696 24812
rect 7380 24828 7432 24880
rect 7840 24828 7892 24880
rect 5264 24624 5316 24676
rect 5632 24624 5684 24676
rect 7012 24735 7064 24744
rect 7012 24701 7021 24735
rect 7021 24701 7055 24735
rect 7055 24701 7064 24735
rect 7012 24692 7064 24701
rect 8668 24828 8720 24880
rect 9588 24828 9640 24880
rect 15936 24828 15988 24880
rect 10048 24803 10100 24812
rect 10048 24769 10057 24803
rect 10057 24769 10091 24803
rect 10091 24769 10100 24803
rect 10048 24760 10100 24769
rect 10508 24760 10560 24812
rect 8668 24692 8720 24744
rect 12256 24692 12308 24744
rect 14648 24803 14700 24812
rect 14648 24769 14657 24803
rect 14657 24769 14691 24803
rect 14691 24769 14700 24803
rect 14648 24760 14700 24769
rect 14740 24760 14792 24812
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 15568 24803 15620 24812
rect 15568 24769 15577 24803
rect 15577 24769 15611 24803
rect 15611 24769 15620 24803
rect 17960 24828 18012 24880
rect 15568 24760 15620 24769
rect 16948 24803 17000 24812
rect 16948 24769 16957 24803
rect 16957 24769 16991 24803
rect 16991 24769 17000 24803
rect 16948 24760 17000 24769
rect 17132 24760 17184 24812
rect 17316 24803 17368 24812
rect 17316 24769 17325 24803
rect 17325 24769 17359 24803
rect 17359 24769 17368 24803
rect 17316 24760 17368 24769
rect 17500 24803 17552 24812
rect 17500 24769 17509 24803
rect 17509 24769 17543 24803
rect 17543 24769 17552 24803
rect 17500 24760 17552 24769
rect 17776 24760 17828 24812
rect 21272 24896 21324 24948
rect 18420 24760 18472 24812
rect 18880 24803 18932 24812
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 18972 24803 19024 24812
rect 18972 24769 18981 24803
rect 18981 24769 19015 24803
rect 19015 24769 19024 24803
rect 18972 24760 19024 24769
rect 19524 24760 19576 24812
rect 20076 24828 20128 24880
rect 22560 24828 22612 24880
rect 23756 24828 23808 24880
rect 24032 24871 24084 24880
rect 24032 24837 24041 24871
rect 24041 24837 24075 24871
rect 24075 24837 24084 24871
rect 24032 24828 24084 24837
rect 25136 24828 25188 24880
rect 27528 24828 27580 24880
rect 19984 24760 20036 24812
rect 21732 24760 21784 24812
rect 2412 24556 2464 24608
rect 6092 24556 6144 24608
rect 7564 24624 7616 24676
rect 7656 24624 7708 24676
rect 8944 24556 8996 24608
rect 9956 24599 10008 24608
rect 9956 24565 9965 24599
rect 9965 24565 9999 24599
rect 9999 24565 10008 24599
rect 9956 24556 10008 24565
rect 10232 24624 10284 24676
rect 11152 24556 11204 24608
rect 11980 24556 12032 24608
rect 14556 24556 14608 24608
rect 14740 24599 14792 24608
rect 14740 24565 14749 24599
rect 14749 24565 14783 24599
rect 14783 24565 14792 24599
rect 14740 24556 14792 24565
rect 15476 24624 15528 24676
rect 16948 24624 17000 24676
rect 17316 24624 17368 24676
rect 17500 24624 17552 24676
rect 19156 24624 19208 24676
rect 19708 24624 19760 24676
rect 16580 24556 16632 24608
rect 17592 24556 17644 24608
rect 17684 24599 17736 24608
rect 17684 24565 17693 24599
rect 17693 24565 17727 24599
rect 17727 24565 17736 24599
rect 17684 24556 17736 24565
rect 19616 24556 19668 24608
rect 22836 24692 22888 24744
rect 20076 24624 20128 24676
rect 20628 24624 20680 24676
rect 21824 24624 21876 24676
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 26240 24803 26292 24812
rect 26240 24769 26249 24803
rect 26249 24769 26283 24803
rect 26283 24769 26292 24803
rect 26240 24760 26292 24769
rect 27160 24760 27212 24812
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 27620 24760 27672 24812
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29276 24760 29328 24769
rect 24216 24692 24268 24744
rect 23664 24599 23716 24608
rect 23664 24565 23673 24599
rect 23673 24565 23707 24599
rect 23707 24565 23716 24599
rect 23664 24556 23716 24565
rect 26332 24599 26384 24608
rect 26332 24565 26341 24599
rect 26341 24565 26375 24599
rect 26375 24565 26384 24599
rect 26332 24556 26384 24565
rect 26792 24556 26844 24608
rect 27804 24624 27856 24676
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 5356 24395 5408 24404
rect 5356 24361 5365 24395
rect 5365 24361 5399 24395
rect 5399 24361 5408 24395
rect 5356 24352 5408 24361
rect 5540 24352 5592 24404
rect 6276 24352 6328 24404
rect 7564 24395 7616 24404
rect 7564 24361 7573 24395
rect 7573 24361 7607 24395
rect 7607 24361 7616 24395
rect 7564 24352 7616 24361
rect 4252 24284 4304 24336
rect 4804 24284 4856 24336
rect 5172 24284 5224 24336
rect 2780 24216 2832 24268
rect 3700 24216 3752 24268
rect 4160 24216 4212 24268
rect 4620 24216 4672 24268
rect 3240 24148 3292 24200
rect 4528 24148 4580 24200
rect 6184 24216 6236 24268
rect 5540 24148 5592 24200
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 6736 24284 6788 24336
rect 7840 24352 7892 24404
rect 8208 24352 8260 24404
rect 6184 24123 6236 24132
rect 3884 24012 3936 24064
rect 4344 24012 4396 24064
rect 6184 24089 6193 24123
rect 6193 24089 6227 24123
rect 6227 24089 6236 24123
rect 6184 24080 6236 24089
rect 6000 24012 6052 24064
rect 7748 24191 7800 24200
rect 7748 24157 7757 24191
rect 7757 24157 7791 24191
rect 7791 24157 7800 24191
rect 7748 24148 7800 24157
rect 8208 24216 8260 24268
rect 8116 24191 8168 24200
rect 8116 24157 8125 24191
rect 8125 24157 8159 24191
rect 8159 24157 8168 24191
rect 8116 24148 8168 24157
rect 9956 24352 10008 24404
rect 13912 24352 13964 24404
rect 8760 24284 8812 24336
rect 14464 24284 14516 24336
rect 14924 24352 14976 24404
rect 16856 24352 16908 24404
rect 16948 24352 17000 24404
rect 17408 24395 17460 24404
rect 17408 24361 17417 24395
rect 17417 24361 17451 24395
rect 17451 24361 17460 24395
rect 17408 24352 17460 24361
rect 17592 24352 17644 24404
rect 18236 24352 18288 24404
rect 8852 24216 8904 24268
rect 8668 24148 8720 24200
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 7932 24123 7984 24132
rect 7932 24089 7941 24123
rect 7941 24089 7975 24123
rect 7975 24089 7984 24123
rect 7932 24080 7984 24089
rect 9772 24148 9824 24200
rect 10232 24216 10284 24268
rect 9956 24191 10008 24200
rect 9956 24157 9965 24191
rect 9965 24157 9999 24191
rect 9999 24157 10008 24191
rect 9956 24148 10008 24157
rect 10416 24216 10468 24268
rect 11980 24191 12032 24200
rect 11980 24157 11990 24191
rect 11990 24157 12024 24191
rect 12024 24157 12032 24191
rect 11980 24148 12032 24157
rect 12164 24191 12216 24200
rect 12164 24157 12173 24191
rect 12173 24157 12207 24191
rect 12207 24157 12216 24191
rect 12164 24148 12216 24157
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 9956 24012 10008 24064
rect 10048 24012 10100 24064
rect 10508 24123 10560 24132
rect 10508 24089 10517 24123
rect 10517 24089 10551 24123
rect 10551 24089 10560 24123
rect 10508 24080 10560 24089
rect 10600 24123 10652 24132
rect 10600 24089 10609 24123
rect 10609 24089 10643 24123
rect 10643 24089 10652 24123
rect 10600 24080 10652 24089
rect 11612 24080 11664 24132
rect 12532 24148 12584 24200
rect 10232 24055 10284 24064
rect 10232 24021 10241 24055
rect 10241 24021 10275 24055
rect 10275 24021 10284 24055
rect 10232 24012 10284 24021
rect 10784 24012 10836 24064
rect 12440 24012 12492 24064
rect 13912 24216 13964 24268
rect 14096 24259 14148 24268
rect 14096 24225 14105 24259
rect 14105 24225 14139 24259
rect 14139 24225 14148 24259
rect 14096 24216 14148 24225
rect 15016 24284 15068 24336
rect 18420 24284 18472 24336
rect 19340 24352 19392 24404
rect 12900 24123 12952 24132
rect 12900 24089 12909 24123
rect 12909 24089 12943 24123
rect 12943 24089 12952 24123
rect 12900 24080 12952 24089
rect 12992 24123 13044 24132
rect 12992 24089 13001 24123
rect 13001 24089 13035 24123
rect 13035 24089 13044 24123
rect 12992 24080 13044 24089
rect 13268 24148 13320 24200
rect 13544 24080 13596 24132
rect 14004 24080 14056 24132
rect 15016 24191 15068 24200
rect 15016 24157 15025 24191
rect 15025 24157 15059 24191
rect 15059 24157 15068 24191
rect 15016 24148 15068 24157
rect 15292 24191 15344 24200
rect 15292 24157 15301 24191
rect 15301 24157 15335 24191
rect 15335 24157 15344 24191
rect 15292 24148 15344 24157
rect 15568 24148 15620 24200
rect 15660 24191 15712 24200
rect 15660 24157 15669 24191
rect 15669 24157 15703 24191
rect 15703 24157 15712 24191
rect 15660 24148 15712 24157
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 16948 24191 17000 24200
rect 16948 24157 16957 24191
rect 16957 24157 16991 24191
rect 16991 24157 17000 24191
rect 16948 24148 17000 24157
rect 17224 24191 17276 24200
rect 17224 24157 17247 24191
rect 17247 24157 17276 24191
rect 17224 24148 17276 24157
rect 14832 24080 14884 24132
rect 13084 24012 13136 24064
rect 13268 24012 13320 24064
rect 13728 24012 13780 24064
rect 17040 24123 17092 24132
rect 17040 24089 17049 24123
rect 17049 24089 17083 24123
rect 17083 24089 17092 24123
rect 17040 24080 17092 24089
rect 17408 24148 17460 24200
rect 17592 24148 17644 24200
rect 18052 24191 18104 24200
rect 18052 24157 18061 24191
rect 18061 24157 18095 24191
rect 18095 24157 18104 24191
rect 18052 24148 18104 24157
rect 18420 24191 18472 24200
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 19340 24216 19392 24268
rect 19984 24284 20036 24336
rect 21088 24284 21140 24336
rect 19708 24148 19760 24200
rect 19248 24080 19300 24132
rect 20536 24191 20588 24194
rect 20536 24157 20545 24191
rect 20545 24157 20579 24191
rect 20579 24157 20588 24191
rect 20536 24142 20588 24157
rect 20076 24080 20128 24132
rect 16672 24055 16724 24064
rect 16672 24021 16681 24055
rect 16681 24021 16715 24055
rect 16715 24021 16724 24055
rect 16672 24012 16724 24021
rect 16948 24012 17000 24064
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 19708 24012 19760 24064
rect 19892 24012 19944 24064
rect 21364 24191 21416 24200
rect 21364 24157 21373 24191
rect 21373 24157 21407 24191
rect 21407 24157 21416 24191
rect 21364 24148 21416 24157
rect 21088 24080 21140 24132
rect 21272 24123 21324 24132
rect 21272 24089 21281 24123
rect 21281 24089 21315 24123
rect 21315 24089 21324 24123
rect 22560 24352 22612 24404
rect 22836 24352 22888 24404
rect 24216 24395 24268 24404
rect 24216 24361 24225 24395
rect 24225 24361 24259 24395
rect 24259 24361 24268 24395
rect 24216 24352 24268 24361
rect 25136 24352 25188 24404
rect 21824 24284 21876 24336
rect 22008 24284 22060 24336
rect 21824 24191 21876 24200
rect 21824 24157 21833 24191
rect 21833 24157 21867 24191
rect 21867 24157 21876 24191
rect 21824 24148 21876 24157
rect 21916 24191 21968 24200
rect 21916 24157 21925 24191
rect 21925 24157 21959 24191
rect 21959 24157 21968 24191
rect 21916 24148 21968 24157
rect 22100 24259 22152 24268
rect 22100 24225 22109 24259
rect 22109 24225 22143 24259
rect 22143 24225 22152 24259
rect 22100 24216 22152 24225
rect 23112 24327 23164 24336
rect 23112 24293 23121 24327
rect 23121 24293 23155 24327
rect 23155 24293 23164 24327
rect 23112 24284 23164 24293
rect 26240 24352 26292 24404
rect 27436 24352 27488 24404
rect 23756 24259 23808 24268
rect 23756 24225 23765 24259
rect 23765 24225 23799 24259
rect 23799 24225 23808 24259
rect 23756 24216 23808 24225
rect 24032 24148 24084 24200
rect 27620 24191 27672 24200
rect 27620 24157 27629 24191
rect 27629 24157 27663 24191
rect 27663 24157 27672 24191
rect 27620 24148 27672 24157
rect 21272 24080 21324 24089
rect 20904 24055 20956 24064
rect 20904 24021 20913 24055
rect 20913 24021 20947 24055
rect 20947 24021 20956 24055
rect 20904 24012 20956 24021
rect 21548 24055 21600 24064
rect 21548 24021 21557 24055
rect 21557 24021 21591 24055
rect 21591 24021 21600 24055
rect 21548 24012 21600 24021
rect 21916 24012 21968 24064
rect 23664 24080 23716 24132
rect 23940 24080 23992 24132
rect 25688 24123 25740 24132
rect 25688 24089 25697 24123
rect 25697 24089 25731 24123
rect 25731 24089 25740 24123
rect 25688 24080 25740 24089
rect 26332 24080 26384 24132
rect 28172 24080 28224 24132
rect 28908 24080 28960 24132
rect 26516 24012 26568 24064
rect 27528 24012 27580 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 3240 23851 3292 23860
rect 3240 23817 3249 23851
rect 3249 23817 3283 23851
rect 3283 23817 3292 23851
rect 3240 23808 3292 23817
rect 4252 23851 4304 23860
rect 4252 23817 4261 23851
rect 4261 23817 4295 23851
rect 4295 23817 4304 23851
rect 4252 23808 4304 23817
rect 4804 23808 4856 23860
rect 7656 23808 7708 23860
rect 8024 23808 8076 23860
rect 4528 23740 4580 23792
rect 848 23672 900 23724
rect 3976 23672 4028 23724
rect 4160 23715 4212 23724
rect 4160 23681 4169 23715
rect 4169 23681 4203 23715
rect 4203 23681 4212 23715
rect 4160 23672 4212 23681
rect 4344 23715 4396 23724
rect 4344 23681 4353 23715
rect 4353 23681 4387 23715
rect 4387 23681 4396 23715
rect 4344 23672 4396 23681
rect 5264 23740 5316 23792
rect 4896 23672 4948 23724
rect 6092 23672 6144 23724
rect 6276 23672 6328 23724
rect 6552 23672 6604 23724
rect 7196 23715 7248 23724
rect 7196 23681 7205 23715
rect 7205 23681 7239 23715
rect 7239 23681 7248 23715
rect 7196 23672 7248 23681
rect 5356 23604 5408 23656
rect 6368 23604 6420 23656
rect 7564 23672 7616 23724
rect 8024 23672 8076 23724
rect 8576 23715 8628 23724
rect 8576 23681 8585 23715
rect 8585 23681 8619 23715
rect 8619 23681 8628 23715
rect 8576 23672 8628 23681
rect 8668 23715 8720 23724
rect 8668 23681 8677 23715
rect 8677 23681 8711 23715
rect 8711 23681 8720 23715
rect 8668 23672 8720 23681
rect 9404 23672 9456 23724
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 9680 23715 9732 23724
rect 9680 23681 9689 23715
rect 9689 23681 9723 23715
rect 9723 23681 9732 23715
rect 9680 23672 9732 23681
rect 9772 23672 9824 23724
rect 11152 23783 11204 23792
rect 11152 23749 11161 23783
rect 11161 23749 11195 23783
rect 11195 23749 11204 23783
rect 11152 23740 11204 23749
rect 10784 23715 10836 23724
rect 4712 23468 4764 23520
rect 6000 23511 6052 23520
rect 6000 23477 6009 23511
rect 6009 23477 6043 23511
rect 6043 23477 6052 23511
rect 6000 23468 6052 23477
rect 6828 23468 6880 23520
rect 7380 23536 7432 23588
rect 8300 23536 8352 23588
rect 8576 23536 8628 23588
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 12532 23740 12584 23792
rect 17960 23808 18012 23860
rect 19248 23808 19300 23860
rect 19524 23808 19576 23860
rect 19708 23851 19760 23860
rect 19708 23817 19717 23851
rect 19717 23817 19751 23851
rect 19751 23817 19760 23851
rect 19708 23808 19760 23817
rect 25688 23808 25740 23860
rect 28172 23851 28224 23860
rect 28172 23817 28181 23851
rect 28181 23817 28215 23851
rect 28215 23817 28224 23851
rect 28172 23808 28224 23817
rect 28908 23851 28960 23860
rect 28908 23817 28917 23851
rect 28917 23817 28951 23851
rect 28951 23817 28960 23851
rect 28908 23808 28960 23817
rect 10232 23536 10284 23588
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 14188 23783 14240 23792
rect 14188 23749 14197 23783
rect 14197 23749 14231 23783
rect 14231 23749 14240 23783
rect 14188 23740 14240 23749
rect 15844 23740 15896 23792
rect 17224 23740 17276 23792
rect 18144 23740 18196 23792
rect 19892 23783 19944 23792
rect 19892 23749 19901 23783
rect 19901 23749 19935 23783
rect 19935 23749 19944 23783
rect 19892 23740 19944 23749
rect 21364 23740 21416 23792
rect 21824 23740 21876 23792
rect 25228 23740 25280 23792
rect 29276 23783 29328 23792
rect 29276 23749 29285 23783
rect 29285 23749 29319 23783
rect 29319 23749 29328 23783
rect 29276 23740 29328 23749
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 13268 23604 13320 23656
rect 13912 23715 13964 23724
rect 13912 23681 13922 23715
rect 13922 23681 13956 23715
rect 13956 23681 13964 23715
rect 13912 23672 13964 23681
rect 14372 23672 14424 23724
rect 14464 23672 14516 23724
rect 15108 23604 15160 23656
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 17500 23672 17552 23724
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 19984 23672 20036 23724
rect 20904 23672 20956 23724
rect 21180 23672 21232 23724
rect 26792 23715 26844 23724
rect 26792 23681 26801 23715
rect 26801 23681 26835 23715
rect 26835 23681 26844 23715
rect 26792 23672 26844 23681
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 27528 23672 27580 23724
rect 29000 23715 29052 23724
rect 29000 23681 29009 23715
rect 29009 23681 29043 23715
rect 29043 23681 29052 23715
rect 29000 23672 29052 23681
rect 19156 23604 19208 23656
rect 9772 23468 9824 23520
rect 9956 23468 10008 23520
rect 11060 23468 11112 23520
rect 11244 23468 11296 23520
rect 13544 23468 13596 23520
rect 16856 23468 16908 23520
rect 16948 23468 17000 23520
rect 18880 23468 18932 23520
rect 19800 23468 19852 23520
rect 19892 23511 19944 23520
rect 19892 23477 19901 23511
rect 19901 23477 19935 23511
rect 19935 23477 19944 23511
rect 19892 23468 19944 23477
rect 20536 23511 20588 23520
rect 20536 23477 20545 23511
rect 20545 23477 20579 23511
rect 20579 23477 20588 23511
rect 20536 23468 20588 23477
rect 21548 23468 21600 23520
rect 27344 23647 27396 23656
rect 27344 23613 27353 23647
rect 27353 23613 27387 23647
rect 27387 23613 27396 23647
rect 27344 23604 27396 23613
rect 27712 23647 27764 23656
rect 27712 23613 27721 23647
rect 27721 23613 27755 23647
rect 27755 23613 27764 23647
rect 27712 23604 27764 23613
rect 27896 23468 27948 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 4620 23264 4672 23316
rect 5632 23264 5684 23316
rect 11244 23264 11296 23316
rect 12256 23307 12308 23316
rect 12256 23273 12265 23307
rect 12265 23273 12299 23307
rect 12299 23273 12308 23307
rect 12256 23264 12308 23273
rect 12992 23264 13044 23316
rect 7196 23196 7248 23248
rect 9772 23196 9824 23248
rect 10600 23196 10652 23248
rect 4436 23128 4488 23180
rect 9312 23128 9364 23180
rect 10876 23128 10928 23180
rect 12440 23171 12492 23180
rect 12440 23137 12449 23171
rect 12449 23137 12483 23171
rect 12483 23137 12492 23171
rect 12440 23128 12492 23137
rect 13912 23196 13964 23248
rect 14096 23196 14148 23248
rect 4804 23060 4856 23112
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5724 23103 5776 23112
rect 5724 23069 5733 23103
rect 5733 23069 5767 23103
rect 5767 23069 5776 23103
rect 5724 23060 5776 23069
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 7472 23103 7524 23112
rect 7472 23069 7482 23103
rect 7482 23069 7516 23103
rect 7516 23069 7524 23103
rect 7472 23060 7524 23069
rect 8024 23060 8076 23112
rect 10048 23060 10100 23112
rect 10232 23060 10284 23112
rect 11060 23103 11112 23112
rect 11060 23069 11069 23103
rect 11069 23069 11103 23103
rect 11103 23069 11112 23103
rect 11060 23060 11112 23069
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 11244 23060 11296 23112
rect 14372 23171 14424 23180
rect 14372 23137 14381 23171
rect 14381 23137 14415 23171
rect 14415 23137 14424 23171
rect 14372 23128 14424 23137
rect 2688 22992 2740 23044
rect 5264 22992 5316 23044
rect 5540 23035 5592 23044
rect 5540 23001 5549 23035
rect 5549 23001 5583 23035
rect 5583 23001 5592 23035
rect 5540 22992 5592 23001
rect 4896 22924 4948 22976
rect 7656 23035 7708 23044
rect 7656 23001 7665 23035
rect 7665 23001 7699 23035
rect 7699 23001 7708 23035
rect 7656 22992 7708 23001
rect 14096 23103 14148 23112
rect 14096 23069 14105 23103
rect 14105 23069 14139 23103
rect 14139 23069 14148 23103
rect 14096 23060 14148 23069
rect 14280 23060 14332 23112
rect 16672 23264 16724 23316
rect 16948 23264 17000 23316
rect 18328 23264 18380 23316
rect 19156 23264 19208 23316
rect 21732 23307 21784 23316
rect 21732 23273 21741 23307
rect 21741 23273 21775 23307
rect 21775 23273 21784 23307
rect 21732 23264 21784 23273
rect 27712 23264 27764 23316
rect 15200 23196 15252 23248
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15476 23060 15528 23112
rect 16396 23103 16448 23112
rect 16396 23069 16405 23103
rect 16405 23069 16439 23103
rect 16439 23069 16448 23103
rect 16396 23060 16448 23069
rect 16672 23105 16724 23112
rect 16672 23071 16681 23105
rect 16681 23071 16715 23105
rect 16715 23071 16724 23105
rect 16672 23060 16724 23071
rect 14740 23035 14792 23044
rect 14740 23001 14749 23035
rect 14749 23001 14783 23035
rect 14783 23001 14792 23035
rect 14740 22992 14792 23001
rect 16856 23035 16908 23044
rect 16856 23001 16865 23035
rect 16865 23001 16899 23035
rect 16899 23001 16908 23035
rect 16856 22992 16908 23001
rect 16948 22992 17000 23044
rect 15108 22967 15160 22976
rect 15108 22933 15117 22967
rect 15117 22933 15151 22967
rect 15151 22933 15160 22967
rect 15108 22924 15160 22933
rect 16672 22924 16724 22976
rect 17960 23103 18012 23112
rect 17960 23069 17969 23103
rect 17969 23069 18003 23103
rect 18003 23069 18012 23103
rect 17960 23060 18012 23069
rect 18052 23103 18104 23112
rect 18052 23069 18061 23103
rect 18061 23069 18095 23103
rect 18095 23069 18104 23103
rect 18052 23060 18104 23069
rect 18328 23060 18380 23112
rect 18696 23103 18748 23112
rect 18696 23069 18705 23103
rect 18705 23069 18739 23103
rect 18739 23069 18748 23103
rect 18696 23060 18748 23069
rect 19064 23196 19116 23248
rect 23848 23196 23900 23248
rect 23572 23128 23624 23180
rect 19432 23060 19484 23112
rect 21732 23060 21784 23112
rect 28172 23128 28224 23180
rect 23664 22992 23716 23044
rect 26240 23060 26292 23112
rect 27160 23103 27212 23112
rect 27160 23069 27169 23103
rect 27169 23069 27203 23103
rect 27203 23069 27212 23103
rect 27160 23060 27212 23069
rect 27344 23103 27396 23112
rect 27344 23069 27353 23103
rect 27353 23069 27387 23103
rect 27387 23069 27396 23103
rect 27344 23060 27396 23069
rect 25412 22992 25464 23044
rect 27712 22992 27764 23044
rect 20444 22924 20496 22976
rect 21456 22924 21508 22976
rect 21824 22924 21876 22976
rect 22008 22924 22060 22976
rect 25044 22967 25096 22976
rect 25044 22933 25053 22967
rect 25053 22933 25087 22967
rect 25087 22933 25096 22967
rect 25044 22924 25096 22933
rect 27896 22967 27948 22976
rect 27896 22933 27905 22967
rect 27905 22933 27939 22967
rect 27939 22933 27948 22967
rect 27896 22924 27948 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 4436 22720 4488 22772
rect 2688 22584 2740 22636
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 4160 22584 4212 22636
rect 4804 22652 4856 22704
rect 5540 22695 5592 22704
rect 5540 22661 5549 22695
rect 5549 22661 5583 22695
rect 5583 22661 5592 22695
rect 5540 22652 5592 22661
rect 848 22516 900 22568
rect 3056 22559 3108 22568
rect 3056 22525 3065 22559
rect 3065 22525 3099 22559
rect 3099 22525 3108 22559
rect 3056 22516 3108 22525
rect 5724 22627 5776 22636
rect 5724 22593 5733 22627
rect 5733 22593 5767 22627
rect 5767 22593 5776 22627
rect 5724 22584 5776 22593
rect 6736 22652 6788 22704
rect 6920 22652 6972 22704
rect 7656 22695 7708 22704
rect 7656 22661 7665 22695
rect 7665 22661 7699 22695
rect 7699 22661 7708 22695
rect 7656 22652 7708 22661
rect 6368 22627 6420 22636
rect 6368 22593 6377 22627
rect 6377 22593 6411 22627
rect 6411 22593 6420 22627
rect 6368 22584 6420 22593
rect 6552 22516 6604 22568
rect 7748 22627 7800 22636
rect 7748 22593 7757 22627
rect 7757 22593 7791 22627
rect 7791 22593 7800 22627
rect 7748 22584 7800 22593
rect 8024 22720 8076 22772
rect 8208 22720 8260 22772
rect 9680 22720 9732 22772
rect 9956 22720 10008 22772
rect 10876 22720 10928 22772
rect 14740 22720 14792 22772
rect 15476 22720 15528 22772
rect 16396 22720 16448 22772
rect 8116 22584 8168 22636
rect 6184 22448 6236 22500
rect 6920 22448 6972 22500
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 5632 22380 5684 22432
rect 7380 22423 7432 22432
rect 7380 22389 7389 22423
rect 7389 22389 7423 22423
rect 7423 22389 7432 22423
rect 7380 22380 7432 22389
rect 8208 22516 8260 22568
rect 7748 22448 7800 22500
rect 8944 22584 8996 22636
rect 10324 22584 10376 22636
rect 10508 22516 10560 22568
rect 10876 22584 10928 22636
rect 12992 22695 13044 22704
rect 12992 22661 13001 22695
rect 13001 22661 13035 22695
rect 13035 22661 13044 22695
rect 12992 22652 13044 22661
rect 14372 22652 14424 22704
rect 16856 22652 16908 22704
rect 17408 22720 17460 22772
rect 17316 22695 17368 22704
rect 17316 22661 17325 22695
rect 17325 22661 17359 22695
rect 17359 22661 17368 22695
rect 17316 22652 17368 22661
rect 18052 22720 18104 22772
rect 12164 22516 12216 22568
rect 12716 22516 12768 22568
rect 13268 22584 13320 22636
rect 16120 22584 16172 22636
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 17684 22627 17736 22636
rect 17684 22593 17694 22627
rect 17694 22593 17728 22627
rect 17728 22593 17736 22627
rect 17684 22584 17736 22593
rect 13728 22516 13780 22568
rect 17960 22695 18012 22704
rect 17960 22661 17969 22695
rect 17969 22661 18003 22695
rect 18003 22661 18012 22695
rect 17960 22652 18012 22661
rect 18328 22695 18380 22704
rect 18328 22661 18337 22695
rect 18337 22661 18371 22695
rect 18371 22661 18380 22695
rect 18328 22652 18380 22661
rect 17868 22516 17920 22568
rect 18420 22584 18472 22636
rect 19708 22720 19760 22772
rect 19432 22652 19484 22704
rect 20168 22652 20220 22704
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 19708 22584 19760 22636
rect 19800 22627 19852 22636
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 21180 22763 21232 22772
rect 21180 22729 21189 22763
rect 21189 22729 21223 22763
rect 21223 22729 21232 22763
rect 21180 22720 21232 22729
rect 21732 22720 21784 22772
rect 23388 22720 23440 22772
rect 20720 22584 20772 22636
rect 20996 22627 21048 22636
rect 20996 22593 21005 22627
rect 21005 22593 21039 22627
rect 21039 22593 21048 22627
rect 20996 22584 21048 22593
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 21732 22584 21784 22636
rect 25412 22763 25464 22772
rect 25412 22729 25421 22763
rect 25421 22729 25455 22763
rect 25455 22729 25464 22763
rect 25412 22720 25464 22729
rect 27712 22720 27764 22772
rect 23940 22695 23992 22704
rect 23940 22661 23949 22695
rect 23949 22661 23983 22695
rect 23983 22661 23992 22695
rect 23940 22652 23992 22661
rect 27896 22695 27948 22704
rect 27896 22661 27905 22695
rect 27905 22661 27939 22695
rect 27939 22661 27948 22695
rect 27896 22652 27948 22661
rect 28908 22652 28960 22704
rect 25044 22584 25096 22636
rect 26240 22584 26292 22636
rect 19892 22516 19944 22568
rect 20260 22516 20312 22568
rect 20444 22516 20496 22568
rect 27620 22559 27672 22568
rect 27620 22525 27629 22559
rect 27629 22525 27663 22559
rect 27663 22525 27672 22559
rect 27620 22516 27672 22525
rect 13544 22448 13596 22500
rect 14740 22448 14792 22500
rect 14924 22448 14976 22500
rect 15384 22448 15436 22500
rect 18696 22448 18748 22500
rect 18880 22448 18932 22500
rect 10784 22380 10836 22432
rect 11704 22423 11756 22432
rect 11704 22389 11713 22423
rect 11713 22389 11747 22423
rect 11747 22389 11756 22423
rect 11704 22380 11756 22389
rect 12532 22380 12584 22432
rect 12900 22380 12952 22432
rect 19064 22380 19116 22432
rect 20536 22423 20588 22432
rect 20536 22389 20545 22423
rect 20545 22389 20579 22423
rect 20579 22389 20588 22423
rect 20536 22380 20588 22389
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 24400 22380 24452 22432
rect 26700 22380 26752 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 3056 22176 3108 22228
rect 4620 22176 4672 22228
rect 5264 22176 5316 22228
rect 2964 22108 3016 22160
rect 6552 22108 6604 22160
rect 4068 22040 4120 22092
rect 6828 22040 6880 22092
rect 7196 22108 7248 22160
rect 7472 22040 7524 22092
rect 7656 22083 7708 22092
rect 7656 22049 7665 22083
rect 7665 22049 7699 22083
rect 7699 22049 7708 22083
rect 7656 22040 7708 22049
rect 4068 21904 4120 21956
rect 3884 21836 3936 21888
rect 5356 21904 5408 21956
rect 4712 21836 4764 21888
rect 6552 21836 6604 21888
rect 6736 22015 6788 22024
rect 6736 21981 6745 22015
rect 6745 21981 6779 22015
rect 6779 21981 6788 22015
rect 6736 21972 6788 21981
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 6828 21947 6880 21956
rect 6828 21913 6837 21947
rect 6837 21913 6871 21947
rect 6871 21913 6880 21947
rect 6828 21904 6880 21913
rect 7288 21904 7340 21956
rect 8208 22040 8260 22092
rect 8484 22040 8536 22092
rect 8668 22040 8720 22092
rect 7104 21879 7156 21888
rect 7104 21845 7113 21879
rect 7113 21845 7147 21879
rect 7147 21845 7156 21879
rect 7104 21836 7156 21845
rect 7932 21836 7984 21888
rect 8300 21972 8352 22024
rect 8392 21947 8444 21956
rect 8392 21913 8401 21947
rect 8401 21913 8435 21947
rect 8435 21913 8444 21947
rect 8392 21904 8444 21913
rect 9312 22083 9364 22092
rect 9312 22049 9321 22083
rect 9321 22049 9355 22083
rect 9355 22049 9364 22083
rect 9312 22040 9364 22049
rect 9772 22040 9824 22092
rect 9128 22015 9180 22024
rect 9128 21981 9137 22015
rect 9137 21981 9171 22015
rect 9171 21981 9180 22015
rect 9128 21972 9180 21981
rect 9404 21904 9456 21956
rect 9588 21836 9640 21888
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 10232 22108 10284 22160
rect 11704 22108 11756 22160
rect 12716 22176 12768 22228
rect 10508 22040 10560 22092
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 10324 21972 10376 21981
rect 10600 21972 10652 22024
rect 10968 21972 11020 22024
rect 11244 22015 11296 22024
rect 11244 21981 11253 22015
rect 11253 21981 11287 22015
rect 11287 21981 11296 22015
rect 11244 21972 11296 21981
rect 12900 22108 12952 22160
rect 13544 22108 13596 22160
rect 14280 22151 14332 22160
rect 14280 22117 14289 22151
rect 14289 22117 14323 22151
rect 14323 22117 14332 22151
rect 14280 22108 14332 22117
rect 15200 22176 15252 22228
rect 17316 22176 17368 22228
rect 19984 22176 20036 22228
rect 20536 22176 20588 22228
rect 11612 21972 11664 22024
rect 12072 21972 12124 22024
rect 12532 22015 12584 22024
rect 13360 22083 13412 22092
rect 13360 22049 13369 22083
rect 13369 22049 13403 22083
rect 13403 22049 13412 22083
rect 13360 22040 13412 22049
rect 11428 21904 11480 21956
rect 11888 21947 11940 21956
rect 11888 21913 11897 21947
rect 11897 21913 11931 21947
rect 11931 21913 11940 21947
rect 11888 21904 11940 21913
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 11980 21904 12032 21913
rect 12532 21981 12571 22015
rect 12571 21981 12584 22015
rect 12532 21972 12584 21981
rect 12440 21904 12492 21956
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 13268 21972 13320 22024
rect 14832 22040 14884 22092
rect 13728 22015 13780 22024
rect 13728 21981 13737 22015
rect 13737 21981 13771 22015
rect 13771 21981 13780 22015
rect 13728 21972 13780 21981
rect 14188 22015 14240 22024
rect 14188 21981 14197 22015
rect 14197 21981 14231 22015
rect 14231 21981 14240 22015
rect 14188 21972 14240 21981
rect 14464 21972 14516 22024
rect 10324 21836 10376 21888
rect 11244 21836 11296 21888
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 11612 21879 11664 21888
rect 11612 21845 11621 21879
rect 11621 21845 11655 21879
rect 11655 21845 11664 21879
rect 11612 21836 11664 21845
rect 11704 21836 11756 21888
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 14924 21972 14976 22024
rect 15384 21972 15436 22024
rect 15660 21972 15712 22024
rect 16764 21972 16816 22024
rect 17132 21972 17184 22024
rect 14832 21904 14884 21956
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 13912 21836 13964 21888
rect 19156 21904 19208 21956
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 17224 21836 17276 21888
rect 17408 21836 17460 21888
rect 19524 22083 19576 22092
rect 19524 22049 19533 22083
rect 19533 22049 19567 22083
rect 19567 22049 19576 22083
rect 19524 22040 19576 22049
rect 19340 21972 19392 22024
rect 19340 21836 19392 21888
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 20720 22108 20772 22160
rect 23848 22176 23900 22228
rect 27160 22176 27212 22228
rect 23388 22108 23440 22160
rect 21732 22040 21784 22092
rect 21824 22040 21876 22092
rect 22560 22040 22612 22092
rect 20076 22015 20128 22024
rect 20076 21981 20085 22015
rect 20085 21981 20119 22015
rect 20119 21981 20128 22015
rect 20076 21972 20128 21981
rect 20260 21972 20312 22024
rect 24492 22083 24544 22092
rect 24492 22049 24501 22083
rect 24501 22049 24535 22083
rect 24535 22049 24544 22083
rect 24492 22040 24544 22049
rect 26056 22040 26108 22092
rect 19892 21947 19944 21956
rect 19892 21913 19901 21947
rect 19901 21913 19935 21947
rect 19935 21913 19944 21947
rect 19892 21904 19944 21913
rect 20168 21904 20220 21956
rect 23572 21947 23624 21956
rect 23572 21913 23581 21947
rect 23581 21913 23615 21947
rect 23615 21913 23624 21947
rect 23572 21904 23624 21913
rect 20628 21836 20680 21888
rect 22928 21836 22980 21888
rect 23112 21879 23164 21888
rect 23112 21845 23121 21879
rect 23121 21845 23155 21879
rect 23155 21845 23164 21879
rect 23112 21836 23164 21845
rect 26608 21972 26660 22024
rect 28908 22083 28960 22092
rect 28908 22049 28917 22083
rect 28917 22049 28951 22083
rect 28951 22049 28960 22083
rect 28908 22040 28960 22049
rect 29000 22015 29052 22024
rect 29000 21981 29009 22015
rect 29009 21981 29043 22015
rect 29043 21981 29052 22015
rect 29000 21972 29052 21981
rect 29276 22015 29328 22024
rect 29276 21981 29285 22015
rect 29285 21981 29319 22015
rect 29319 21981 29328 22015
rect 29276 21972 29328 21981
rect 26700 21904 26752 21956
rect 27068 21836 27120 21888
rect 27160 21879 27212 21888
rect 27160 21845 27169 21879
rect 27169 21845 27203 21879
rect 27203 21845 27212 21879
rect 27160 21836 27212 21845
rect 29184 21879 29236 21888
rect 29184 21845 29193 21879
rect 29193 21845 29227 21879
rect 29227 21845 29236 21879
rect 29184 21836 29236 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 3884 21564 3936 21616
rect 848 21496 900 21548
rect 2780 21496 2832 21548
rect 5540 21496 5592 21548
rect 6644 21632 6696 21684
rect 6000 21564 6052 21616
rect 6460 21496 6512 21548
rect 6644 21539 6696 21548
rect 6644 21505 6653 21539
rect 6653 21505 6687 21539
rect 6687 21505 6696 21539
rect 6644 21496 6696 21505
rect 7932 21632 7984 21684
rect 8392 21632 8444 21684
rect 3148 21471 3200 21480
rect 3148 21437 3157 21471
rect 3157 21437 3191 21471
rect 3191 21437 3200 21471
rect 3148 21428 3200 21437
rect 4620 21428 4672 21480
rect 7196 21428 7248 21480
rect 1768 21360 1820 21412
rect 6552 21360 6604 21412
rect 6644 21360 6696 21412
rect 8484 21564 8536 21616
rect 10232 21632 10284 21684
rect 10600 21632 10652 21684
rect 11612 21632 11664 21684
rect 15292 21632 15344 21684
rect 15568 21632 15620 21684
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 8576 21496 8628 21548
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9588 21539 9640 21548
rect 9588 21505 9597 21539
rect 9597 21505 9631 21539
rect 9631 21505 9640 21539
rect 9588 21496 9640 21505
rect 10600 21496 10652 21548
rect 13452 21564 13504 21616
rect 14280 21564 14332 21616
rect 9956 21428 10008 21480
rect 11612 21496 11664 21548
rect 11980 21496 12032 21548
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 12532 21428 12584 21480
rect 12624 21428 12676 21480
rect 13268 21496 13320 21548
rect 13728 21428 13780 21480
rect 14556 21539 14608 21548
rect 14556 21505 14565 21539
rect 14565 21505 14599 21539
rect 14599 21505 14608 21539
rect 14556 21496 14608 21505
rect 14740 21496 14792 21548
rect 15200 21496 15252 21548
rect 15476 21496 15528 21548
rect 15568 21471 15620 21480
rect 15568 21437 15577 21471
rect 15577 21437 15611 21471
rect 15611 21437 15620 21471
rect 15568 21428 15620 21437
rect 16396 21564 16448 21616
rect 21088 21632 21140 21684
rect 22100 21632 22152 21684
rect 24492 21632 24544 21684
rect 26240 21632 26292 21684
rect 27160 21632 27212 21684
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17316 21539 17368 21548
rect 17316 21505 17325 21539
rect 17325 21505 17359 21539
rect 17359 21505 17368 21539
rect 17316 21496 17368 21505
rect 17684 21496 17736 21548
rect 18788 21539 18840 21548
rect 18788 21505 18797 21539
rect 18797 21505 18831 21539
rect 18831 21505 18840 21539
rect 18788 21496 18840 21505
rect 20996 21564 21048 21616
rect 26332 21564 26384 21616
rect 28816 21564 28868 21616
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 19524 21496 19576 21548
rect 20904 21496 20956 21548
rect 21824 21539 21876 21548
rect 21824 21505 21833 21539
rect 21833 21505 21867 21539
rect 21867 21505 21876 21539
rect 21824 21496 21876 21505
rect 22928 21539 22980 21548
rect 22928 21505 22937 21539
rect 22937 21505 22971 21539
rect 22971 21505 22980 21539
rect 22928 21496 22980 21505
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 23204 21539 23256 21548
rect 23204 21505 23213 21539
rect 23213 21505 23247 21539
rect 23247 21505 23256 21539
rect 23204 21496 23256 21505
rect 23480 21496 23532 21548
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 24216 21496 24268 21548
rect 9128 21360 9180 21412
rect 11244 21360 11296 21412
rect 13268 21360 13320 21412
rect 17040 21360 17092 21412
rect 19984 21428 20036 21480
rect 20812 21360 20864 21412
rect 26240 21539 26292 21548
rect 26240 21505 26249 21539
rect 26249 21505 26283 21539
rect 26283 21505 26292 21539
rect 26240 21496 26292 21505
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 26056 21360 26108 21412
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27528 21539 27580 21548
rect 27528 21505 27537 21539
rect 27537 21505 27571 21539
rect 27571 21505 27580 21539
rect 27528 21496 27580 21505
rect 27344 21403 27396 21412
rect 27344 21369 27353 21403
rect 27353 21369 27387 21403
rect 27387 21369 27396 21403
rect 27344 21360 27396 21369
rect 6828 21292 6880 21344
rect 7380 21292 7432 21344
rect 8668 21292 8720 21344
rect 10508 21292 10560 21344
rect 11888 21292 11940 21344
rect 13360 21292 13412 21344
rect 14464 21292 14516 21344
rect 16304 21292 16356 21344
rect 16580 21292 16632 21344
rect 17132 21335 17184 21344
rect 17132 21301 17141 21335
rect 17141 21301 17175 21335
rect 17175 21301 17184 21335
rect 17132 21292 17184 21301
rect 17316 21292 17368 21344
rect 19064 21292 19116 21344
rect 19616 21292 19668 21344
rect 23756 21292 23808 21344
rect 25320 21292 25372 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 3884 21088 3936 21140
rect 6276 21088 6328 21140
rect 6736 21088 6788 21140
rect 7472 21088 7524 21140
rect 8668 21088 8720 21140
rect 9312 21088 9364 21140
rect 9956 21131 10008 21140
rect 9956 21097 9965 21131
rect 9965 21097 9999 21131
rect 9999 21097 10008 21131
rect 9956 21088 10008 21097
rect 5816 20952 5868 21004
rect 6184 20952 6236 21004
rect 6920 20952 6972 21004
rect 8208 20952 8260 21004
rect 4068 20884 4120 20936
rect 6092 20927 6144 20936
rect 6092 20893 6096 20927
rect 6096 20893 6130 20927
rect 6130 20893 6144 20927
rect 6092 20884 6144 20893
rect 6460 20927 6512 20936
rect 6460 20893 6468 20927
rect 6468 20893 6502 20927
rect 6502 20893 6512 20927
rect 6460 20884 6512 20893
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 6828 20927 6880 20936
rect 6828 20893 6837 20927
rect 6837 20893 6871 20927
rect 6871 20893 6880 20927
rect 6828 20884 6880 20893
rect 7288 20884 7340 20936
rect 8392 20884 8444 20936
rect 9220 20927 9272 20936
rect 9220 20893 9229 20927
rect 9229 20893 9263 20927
rect 9263 20893 9272 20927
rect 9220 20884 9272 20893
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 9496 20884 9548 20936
rect 9956 20884 10008 20936
rect 11520 21020 11572 21072
rect 1400 20816 1452 20868
rect 2780 20816 2832 20868
rect 3516 20816 3568 20868
rect 6184 20859 6236 20868
rect 6184 20825 6193 20859
rect 6193 20825 6227 20859
rect 6227 20825 6236 20859
rect 6184 20816 6236 20825
rect 6368 20816 6420 20868
rect 6920 20859 6972 20868
rect 5908 20791 5960 20800
rect 5908 20757 5917 20791
rect 5917 20757 5951 20791
rect 5951 20757 5960 20791
rect 5908 20748 5960 20757
rect 6000 20748 6052 20800
rect 6920 20825 6929 20859
rect 6929 20825 6963 20859
rect 6963 20825 6972 20859
rect 6920 20816 6972 20825
rect 6552 20748 6604 20800
rect 8944 20816 8996 20868
rect 9680 20859 9732 20868
rect 9680 20825 9689 20859
rect 9689 20825 9723 20859
rect 9723 20825 9732 20859
rect 9680 20816 9732 20825
rect 11888 20927 11940 20936
rect 11888 20893 11897 20927
rect 11897 20893 11931 20927
rect 11931 20893 11940 20927
rect 11888 20884 11940 20893
rect 12992 21088 13044 21140
rect 15568 21088 15620 21140
rect 20352 21088 20404 21140
rect 23204 21131 23256 21140
rect 23204 21097 23213 21131
rect 23213 21097 23247 21131
rect 23247 21097 23256 21131
rect 23204 21088 23256 21097
rect 26424 21088 26476 21140
rect 14372 21020 14424 21072
rect 15476 21020 15528 21072
rect 18788 21020 18840 21072
rect 16488 20952 16540 21004
rect 17224 20952 17276 21004
rect 12808 20927 12860 20936
rect 12808 20893 12817 20927
rect 12817 20893 12851 20927
rect 12851 20893 12860 20927
rect 12808 20884 12860 20893
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 17040 20927 17092 20936
rect 17040 20893 17049 20927
rect 17049 20893 17083 20927
rect 17083 20893 17092 20927
rect 17040 20884 17092 20893
rect 17960 20927 18012 20936
rect 17960 20893 17969 20927
rect 17969 20893 18003 20927
rect 18003 20893 18012 20927
rect 17960 20884 18012 20893
rect 18052 20927 18104 20936
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 10968 20816 11020 20868
rect 11336 20816 11388 20868
rect 11796 20859 11848 20868
rect 11796 20825 11805 20859
rect 11805 20825 11839 20859
rect 11839 20825 11848 20859
rect 11796 20816 11848 20825
rect 16212 20816 16264 20868
rect 18236 20859 18288 20868
rect 18236 20825 18245 20859
rect 18245 20825 18279 20859
rect 18279 20825 18288 20859
rect 18236 20816 18288 20825
rect 19064 20952 19116 21004
rect 21088 21020 21140 21072
rect 23572 21063 23624 21072
rect 23572 21029 23581 21063
rect 23581 21029 23615 21063
rect 23615 21029 23624 21063
rect 23572 21020 23624 21029
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 19524 20884 19576 20936
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 20628 20859 20680 20868
rect 20628 20825 20637 20859
rect 20637 20825 20671 20859
rect 20671 20825 20680 20859
rect 20628 20816 20680 20825
rect 11888 20748 11940 20800
rect 12440 20748 12492 20800
rect 13544 20748 13596 20800
rect 16672 20748 16724 20800
rect 16856 20791 16908 20800
rect 16856 20757 16865 20791
rect 16865 20757 16899 20791
rect 16899 20757 16908 20791
rect 16856 20748 16908 20757
rect 16948 20748 17000 20800
rect 20260 20791 20312 20800
rect 20260 20757 20269 20791
rect 20269 20757 20303 20791
rect 20303 20757 20312 20791
rect 20260 20748 20312 20757
rect 20812 20927 20864 20936
rect 20812 20893 20820 20927
rect 20820 20893 20854 20927
rect 20854 20893 20864 20927
rect 20812 20884 20864 20893
rect 21732 20952 21784 21004
rect 22100 20952 22152 21004
rect 23940 20995 23992 21004
rect 23940 20961 23949 20995
rect 23949 20961 23983 20995
rect 23983 20961 23992 20995
rect 23940 20952 23992 20961
rect 26332 20952 26384 21004
rect 27344 21088 27396 21140
rect 28816 21088 28868 21140
rect 24400 20927 24452 20936
rect 24400 20893 24409 20927
rect 24409 20893 24443 20927
rect 24443 20893 24452 20927
rect 24400 20884 24452 20893
rect 24492 20884 24544 20936
rect 21180 20859 21232 20868
rect 21180 20825 21189 20859
rect 21189 20825 21223 20859
rect 21223 20825 21232 20859
rect 21180 20816 21232 20825
rect 21732 20859 21784 20868
rect 21732 20825 21741 20859
rect 21741 20825 21775 20859
rect 21775 20825 21784 20859
rect 21732 20816 21784 20825
rect 22468 20816 22520 20868
rect 23112 20816 23164 20868
rect 20904 20748 20956 20800
rect 20996 20748 21048 20800
rect 23480 20791 23532 20800
rect 23480 20757 23489 20791
rect 23489 20757 23523 20791
rect 23523 20757 23532 20791
rect 25320 20859 25372 20868
rect 25320 20825 25329 20859
rect 25329 20825 25363 20859
rect 25363 20825 25372 20859
rect 25320 20816 25372 20825
rect 26332 20816 26384 20868
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27160 20816 27212 20868
rect 23480 20748 23532 20757
rect 24860 20748 24912 20800
rect 26056 20748 26108 20800
rect 29000 20884 29052 20936
rect 29276 20927 29328 20936
rect 29276 20893 29285 20927
rect 29285 20893 29319 20927
rect 29319 20893 29328 20927
rect 29276 20884 29328 20893
rect 29828 20748 29880 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 6828 20544 6880 20596
rect 4804 20476 4856 20528
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 5632 20451 5684 20460
rect 5632 20417 5641 20451
rect 5641 20417 5675 20451
rect 5675 20417 5684 20451
rect 5632 20408 5684 20417
rect 7104 20476 7156 20528
rect 6920 20408 6972 20460
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 6184 20340 6236 20392
rect 7196 20340 7248 20392
rect 8116 20408 8168 20460
rect 8576 20476 8628 20528
rect 9312 20544 9364 20596
rect 9496 20544 9548 20596
rect 8944 20451 8996 20460
rect 8944 20417 8951 20451
rect 8951 20417 8996 20451
rect 8944 20408 8996 20417
rect 9128 20451 9180 20460
rect 9128 20417 9137 20451
rect 9137 20417 9171 20451
rect 9171 20417 9180 20451
rect 9128 20408 9180 20417
rect 9220 20451 9272 20460
rect 9680 20476 9732 20528
rect 9220 20417 9234 20451
rect 9234 20417 9268 20451
rect 9268 20417 9272 20451
rect 9220 20408 9272 20417
rect 10784 20544 10836 20596
rect 10048 20476 10100 20528
rect 10692 20476 10744 20528
rect 10232 20408 10284 20460
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 9404 20340 9456 20392
rect 9772 20340 9824 20392
rect 9864 20340 9916 20392
rect 11704 20476 11756 20528
rect 12164 20476 12216 20528
rect 11336 20408 11388 20460
rect 11980 20451 12032 20460
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 5908 20204 5960 20256
rect 6368 20204 6420 20256
rect 7932 20272 7984 20324
rect 8116 20272 8168 20324
rect 8392 20315 8444 20324
rect 8392 20281 8401 20315
rect 8401 20281 8435 20315
rect 8435 20281 8444 20315
rect 8392 20272 8444 20281
rect 9036 20272 9088 20324
rect 9496 20272 9548 20324
rect 12348 20408 12400 20460
rect 13084 20451 13136 20460
rect 13084 20417 13093 20451
rect 13093 20417 13127 20451
rect 13127 20417 13136 20451
rect 13084 20408 13136 20417
rect 13360 20451 13412 20460
rect 13360 20417 13369 20451
rect 13369 20417 13403 20451
rect 13403 20417 13412 20451
rect 13360 20408 13412 20417
rect 13820 20519 13872 20528
rect 13820 20485 13829 20519
rect 13829 20485 13863 20519
rect 13863 20485 13872 20519
rect 13820 20476 13872 20485
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 13636 20408 13688 20460
rect 13912 20451 13964 20460
rect 13912 20417 13921 20451
rect 13921 20417 13955 20451
rect 13955 20417 13964 20451
rect 13912 20408 13964 20417
rect 14188 20451 14240 20460
rect 14188 20417 14197 20451
rect 14197 20417 14231 20451
rect 14231 20417 14240 20451
rect 14188 20408 14240 20417
rect 14556 20544 14608 20596
rect 15016 20476 15068 20528
rect 19432 20544 19484 20596
rect 19984 20544 20036 20596
rect 14556 20451 14608 20460
rect 14556 20417 14566 20451
rect 14566 20417 14600 20451
rect 14600 20417 14608 20451
rect 14556 20408 14608 20417
rect 14924 20451 14976 20460
rect 14924 20417 14938 20451
rect 14938 20417 14972 20451
rect 14972 20417 14976 20451
rect 14924 20408 14976 20417
rect 15108 20408 15160 20460
rect 7840 20204 7892 20256
rect 12348 20272 12400 20324
rect 11520 20204 11572 20256
rect 11704 20204 11756 20256
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17132 20408 17184 20460
rect 14372 20272 14424 20324
rect 16396 20340 16448 20392
rect 17040 20383 17092 20392
rect 17040 20349 17049 20383
rect 17049 20349 17083 20383
rect 17083 20349 17092 20383
rect 17040 20340 17092 20349
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 18328 20408 18380 20460
rect 18696 20408 18748 20460
rect 19340 20451 19392 20460
rect 19340 20417 19349 20451
rect 19349 20417 19383 20451
rect 19383 20417 19392 20451
rect 19340 20408 19392 20417
rect 19524 20451 19576 20460
rect 19524 20417 19534 20451
rect 19534 20417 19568 20451
rect 19568 20417 19576 20451
rect 19524 20408 19576 20417
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 17500 20272 17552 20324
rect 20168 20451 20220 20460
rect 20168 20417 20177 20451
rect 20177 20417 20211 20451
rect 20211 20417 20220 20451
rect 20168 20408 20220 20417
rect 20628 20408 20680 20460
rect 21180 20544 21232 20596
rect 22468 20544 22520 20596
rect 24492 20587 24544 20596
rect 24492 20553 24501 20587
rect 24501 20553 24535 20587
rect 24535 20553 24544 20587
rect 24492 20544 24544 20553
rect 26332 20544 26384 20596
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 21180 20451 21232 20460
rect 21180 20417 21189 20451
rect 21189 20417 21223 20451
rect 21223 20417 21232 20451
rect 21180 20408 21232 20417
rect 21364 20408 21416 20460
rect 22560 20408 22612 20460
rect 29000 20476 29052 20528
rect 19340 20272 19392 20324
rect 19524 20272 19576 20324
rect 16212 20204 16264 20256
rect 16948 20204 17000 20256
rect 17868 20204 17920 20256
rect 19800 20204 19852 20256
rect 20720 20204 20772 20256
rect 21824 20340 21876 20392
rect 22192 20340 22244 20392
rect 27528 20451 27580 20460
rect 27528 20417 27537 20451
rect 27537 20417 27571 20451
rect 27571 20417 27580 20451
rect 27528 20408 27580 20417
rect 22560 20272 22612 20324
rect 24952 20340 25004 20392
rect 27712 20340 27764 20392
rect 29092 20272 29144 20324
rect 27896 20204 27948 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 4804 20000 4856 20052
rect 6184 20043 6236 20052
rect 6184 20009 6193 20043
rect 6193 20009 6227 20043
rect 6227 20009 6236 20043
rect 6184 20000 6236 20009
rect 7932 20000 7984 20052
rect 4896 19932 4948 19984
rect 6460 19932 6512 19984
rect 6736 19932 6788 19984
rect 8944 20000 8996 20052
rect 9864 20000 9916 20052
rect 11244 20000 11296 20052
rect 11520 20000 11572 20052
rect 6644 19907 6696 19916
rect 6644 19873 6653 19907
rect 6653 19873 6687 19907
rect 6687 19873 6696 19907
rect 6644 19864 6696 19873
rect 848 19796 900 19848
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2872 19796 2924 19848
rect 4068 19796 4120 19848
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 6276 19839 6328 19848
rect 6276 19805 6285 19839
rect 6285 19805 6319 19839
rect 6319 19805 6328 19839
rect 6276 19796 6328 19805
rect 6368 19839 6420 19848
rect 6368 19805 6377 19839
rect 6377 19805 6411 19839
rect 6411 19805 6420 19839
rect 6368 19796 6420 19805
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 7472 19907 7524 19916
rect 7472 19873 7481 19907
rect 7481 19873 7515 19907
rect 7515 19873 7524 19907
rect 7472 19864 7524 19873
rect 3424 19728 3476 19780
rect 6460 19728 6512 19780
rect 7288 19796 7340 19848
rect 7840 19864 7892 19916
rect 8116 19796 8168 19848
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 11336 19932 11388 19984
rect 8484 19864 8536 19916
rect 9496 19864 9548 19916
rect 1676 19660 1728 19712
rect 2596 19703 2648 19712
rect 2596 19669 2605 19703
rect 2605 19669 2639 19703
rect 2639 19669 2648 19703
rect 2596 19660 2648 19669
rect 7012 19660 7064 19712
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 8024 19703 8076 19712
rect 8024 19669 8033 19703
rect 8033 19669 8067 19703
rect 8067 19669 8076 19703
rect 8024 19660 8076 19669
rect 8300 19771 8352 19780
rect 8300 19737 8309 19771
rect 8309 19737 8343 19771
rect 8343 19737 8352 19771
rect 8300 19728 8352 19737
rect 9772 19796 9824 19848
rect 10048 19796 10100 19848
rect 9128 19728 9180 19780
rect 9496 19728 9548 19780
rect 9680 19728 9732 19780
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 10784 19839 10836 19848
rect 10784 19805 10793 19839
rect 10793 19805 10827 19839
rect 10827 19805 10836 19839
rect 10784 19796 10836 19805
rect 11704 19907 11756 19916
rect 11704 19873 11713 19907
rect 11713 19873 11747 19907
rect 11747 19873 11756 19907
rect 11704 19864 11756 19873
rect 16672 20000 16724 20052
rect 16764 20000 16816 20052
rect 16948 20000 17000 20052
rect 17316 20000 17368 20052
rect 18144 20000 18196 20052
rect 19432 20000 19484 20052
rect 19892 20000 19944 20052
rect 10600 19728 10652 19780
rect 11244 19796 11296 19848
rect 8760 19660 8812 19712
rect 11980 19728 12032 19780
rect 13360 19796 13412 19848
rect 14740 19932 14792 19984
rect 16212 19932 16264 19984
rect 17132 19932 17184 19984
rect 18052 19932 18104 19984
rect 19800 19975 19852 19984
rect 19800 19941 19809 19975
rect 19809 19941 19843 19975
rect 19843 19941 19852 19975
rect 19800 19932 19852 19941
rect 12992 19660 13044 19712
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 13176 19660 13228 19669
rect 14556 19660 14608 19712
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 21732 20000 21784 20052
rect 21180 19932 21232 19984
rect 21916 19932 21968 19984
rect 14924 19839 14976 19848
rect 14924 19805 14933 19839
rect 14933 19805 14967 19839
rect 14967 19805 14976 19839
rect 14924 19796 14976 19805
rect 15108 19839 15160 19848
rect 15108 19805 15122 19839
rect 15122 19805 15156 19839
rect 15156 19805 15160 19839
rect 15108 19796 15160 19805
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 17408 19796 17460 19848
rect 17592 19796 17644 19848
rect 15016 19771 15068 19780
rect 15016 19737 15025 19771
rect 15025 19737 15059 19771
rect 15059 19737 15068 19771
rect 15016 19728 15068 19737
rect 16672 19728 16724 19780
rect 17500 19728 17552 19780
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18328 19796 18380 19848
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 17960 19728 18012 19780
rect 18236 19728 18288 19780
rect 18788 19771 18840 19780
rect 18788 19737 18797 19771
rect 18797 19737 18831 19771
rect 18831 19737 18840 19771
rect 18788 19728 18840 19737
rect 18972 19839 19024 19848
rect 18972 19805 18981 19839
rect 18981 19805 19015 19839
rect 19015 19805 19024 19839
rect 18972 19796 19024 19805
rect 19616 19839 19668 19848
rect 19616 19805 19637 19839
rect 19637 19805 19668 19839
rect 19616 19796 19668 19805
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 19248 19728 19300 19780
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 22284 19864 22336 19916
rect 23296 19864 23348 19916
rect 26240 19864 26292 19916
rect 26884 19864 26936 19916
rect 27528 20000 27580 20052
rect 27344 19864 27396 19916
rect 21364 19796 21416 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 22836 19796 22888 19848
rect 26976 19839 27028 19848
rect 26976 19805 26985 19839
rect 26985 19805 27019 19839
rect 27019 19805 27028 19839
rect 26976 19796 27028 19805
rect 27620 19907 27672 19916
rect 27620 19873 27629 19907
rect 27629 19873 27663 19907
rect 27663 19873 27672 19907
rect 27620 19864 27672 19873
rect 27896 19907 27948 19916
rect 27896 19873 27905 19907
rect 27905 19873 27939 19907
rect 27939 19873 27948 19907
rect 27896 19864 27948 19873
rect 25136 19728 25188 19780
rect 25964 19728 26016 19780
rect 27252 19728 27304 19780
rect 28908 19728 28960 19780
rect 20812 19660 20864 19712
rect 21640 19703 21692 19712
rect 21640 19669 21649 19703
rect 21649 19669 21683 19703
rect 21683 19669 21692 19703
rect 21640 19660 21692 19669
rect 21824 19660 21876 19712
rect 26792 19703 26844 19712
rect 26792 19669 26801 19703
rect 26801 19669 26835 19703
rect 26835 19669 26844 19703
rect 26792 19660 26844 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 7472 19499 7524 19508
rect 7472 19465 7481 19499
rect 7481 19465 7515 19499
rect 7515 19465 7524 19499
rect 7472 19456 7524 19465
rect 8668 19456 8720 19508
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 10600 19456 10652 19508
rect 10692 19456 10744 19508
rect 1676 19431 1728 19440
rect 1676 19397 1685 19431
rect 1685 19397 1719 19431
rect 1719 19397 1728 19431
rect 1676 19388 1728 19397
rect 3424 19431 3476 19440
rect 3424 19397 3433 19431
rect 3433 19397 3467 19431
rect 3467 19397 3476 19431
rect 3424 19388 3476 19397
rect 5540 19388 5592 19440
rect 8024 19388 8076 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2780 19320 2832 19372
rect 3792 19320 3844 19372
rect 5080 19363 5132 19372
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 6920 19320 6972 19329
rect 7012 19363 7064 19372
rect 7012 19329 7021 19363
rect 7021 19329 7055 19363
rect 7055 19329 7064 19363
rect 7012 19320 7064 19329
rect 7380 19320 7432 19372
rect 4896 19252 4948 19304
rect 7012 19184 7064 19236
rect 7748 19252 7800 19304
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 9128 19388 9180 19440
rect 9864 19431 9916 19440
rect 9864 19397 9873 19431
rect 9873 19397 9907 19431
rect 9907 19397 9916 19431
rect 9864 19388 9916 19397
rect 8668 19320 8720 19372
rect 9404 19320 9456 19372
rect 10508 19320 10560 19372
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 15200 19456 15252 19508
rect 17132 19456 17184 19508
rect 13268 19388 13320 19440
rect 14096 19388 14148 19440
rect 10968 19320 11020 19329
rect 9864 19252 9916 19304
rect 10232 19252 10284 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 12348 19252 12400 19304
rect 12164 19184 12216 19236
rect 13176 19320 13228 19372
rect 14188 19320 14240 19372
rect 17316 19388 17368 19440
rect 14740 19320 14792 19372
rect 15016 19320 15068 19372
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17500 19320 17552 19372
rect 18236 19499 18288 19508
rect 18236 19465 18245 19499
rect 18245 19465 18279 19499
rect 18279 19465 18288 19499
rect 18236 19456 18288 19465
rect 20444 19456 20496 19508
rect 20628 19499 20680 19508
rect 20628 19465 20637 19499
rect 20637 19465 20671 19499
rect 20671 19465 20680 19499
rect 20628 19456 20680 19465
rect 17868 19431 17920 19440
rect 17868 19397 17877 19431
rect 17877 19397 17911 19431
rect 17911 19397 17920 19431
rect 17868 19388 17920 19397
rect 17960 19431 18012 19440
rect 17960 19397 17969 19431
rect 17969 19397 18003 19431
rect 18003 19397 18012 19431
rect 17960 19388 18012 19397
rect 18880 19388 18932 19440
rect 19432 19431 19484 19440
rect 19432 19397 19441 19431
rect 19441 19397 19475 19431
rect 19475 19397 19484 19431
rect 19432 19388 19484 19397
rect 19892 19388 19944 19440
rect 21640 19456 21692 19508
rect 22836 19456 22888 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 25964 19499 26016 19508
rect 25964 19465 25973 19499
rect 25973 19465 26007 19499
rect 26007 19465 26016 19499
rect 25964 19456 26016 19465
rect 27252 19499 27304 19508
rect 27252 19465 27261 19499
rect 27261 19465 27295 19499
rect 27295 19465 27304 19499
rect 27252 19456 27304 19465
rect 27344 19499 27396 19508
rect 27344 19465 27353 19499
rect 27353 19465 27387 19499
rect 27387 19465 27396 19499
rect 27344 19456 27396 19465
rect 27712 19499 27764 19508
rect 27712 19465 27721 19499
rect 27721 19465 27755 19499
rect 27755 19465 27764 19499
rect 27712 19456 27764 19465
rect 28908 19499 28960 19508
rect 28908 19465 28917 19499
rect 28917 19465 28951 19499
rect 28951 19465 28960 19499
rect 28908 19456 28960 19465
rect 21364 19431 21416 19440
rect 21364 19397 21373 19431
rect 21373 19397 21407 19431
rect 21407 19397 21416 19431
rect 21364 19388 21416 19397
rect 18328 19320 18380 19372
rect 18972 19320 19024 19372
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14648 19295 14700 19304
rect 14648 19261 14657 19295
rect 14657 19261 14691 19295
rect 14691 19261 14700 19295
rect 14648 19252 14700 19261
rect 16764 19252 16816 19304
rect 19340 19320 19392 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 19708 19320 19760 19372
rect 20076 19363 20128 19372
rect 20076 19329 20086 19363
rect 20086 19329 20120 19363
rect 20120 19329 20128 19363
rect 20076 19320 20128 19329
rect 14280 19184 14332 19236
rect 16028 19184 16080 19236
rect 16948 19184 17000 19236
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 15292 19116 15344 19168
rect 15844 19116 15896 19168
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 20628 19320 20680 19372
rect 20812 19320 20864 19372
rect 20996 19363 21048 19372
rect 20996 19329 21005 19363
rect 21005 19329 21039 19363
rect 21039 19329 21048 19363
rect 20996 19320 21048 19329
rect 21456 19363 21508 19372
rect 21456 19329 21465 19363
rect 21465 19329 21499 19363
rect 21499 19329 21508 19363
rect 21456 19320 21508 19329
rect 23296 19388 23348 19440
rect 29276 19431 29328 19440
rect 29276 19397 29285 19431
rect 29285 19397 29319 19431
rect 29319 19397 29328 19431
rect 29276 19388 29328 19397
rect 24676 19320 24728 19372
rect 24952 19363 25004 19372
rect 24952 19329 24961 19363
rect 24961 19329 24995 19363
rect 24995 19329 25004 19363
rect 24952 19320 25004 19329
rect 26240 19320 26292 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 22468 19252 22520 19304
rect 26056 19252 26108 19304
rect 29000 19363 29052 19372
rect 29000 19329 29009 19363
rect 29009 19329 29043 19363
rect 29043 19329 29052 19363
rect 29000 19320 29052 19329
rect 26792 19184 26844 19236
rect 26884 19184 26936 19236
rect 27528 19227 27580 19236
rect 27528 19193 27537 19227
rect 27537 19193 27571 19227
rect 27571 19193 27580 19227
rect 27528 19184 27580 19193
rect 21088 19116 21140 19168
rect 29644 19116 29696 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 2780 18912 2832 18964
rect 3148 18912 3200 18964
rect 4344 18912 4396 18964
rect 4896 18912 4948 18964
rect 6460 18912 6512 18964
rect 6920 18912 6972 18964
rect 7196 18955 7248 18964
rect 7196 18921 7205 18955
rect 7205 18921 7239 18955
rect 7239 18921 7248 18955
rect 7196 18912 7248 18921
rect 7288 18912 7340 18964
rect 9496 18912 9548 18964
rect 10508 18955 10560 18964
rect 10508 18921 10517 18955
rect 10517 18921 10551 18955
rect 10551 18921 10560 18955
rect 10508 18912 10560 18921
rect 5080 18887 5132 18896
rect 5080 18853 5089 18887
rect 5089 18853 5123 18887
rect 5123 18853 5132 18887
rect 5080 18844 5132 18853
rect 4160 18776 4212 18828
rect 4252 18776 4304 18828
rect 5724 18844 5776 18896
rect 848 18708 900 18760
rect 2872 18708 2924 18760
rect 4068 18751 4120 18760
rect 4068 18717 4077 18751
rect 4077 18717 4111 18751
rect 4111 18717 4120 18751
rect 4068 18708 4120 18717
rect 4804 18708 4856 18760
rect 5632 18776 5684 18828
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 8668 18844 8720 18896
rect 9680 18844 9732 18896
rect 10968 18844 11020 18896
rect 16856 18912 16908 18964
rect 18144 18912 18196 18964
rect 18696 18912 18748 18964
rect 21088 18912 21140 18964
rect 22468 18955 22520 18964
rect 22468 18921 22477 18955
rect 22477 18921 22511 18955
rect 22511 18921 22520 18955
rect 22468 18912 22520 18921
rect 7104 18708 7156 18760
rect 7288 18751 7340 18760
rect 7288 18717 7297 18751
rect 7297 18717 7331 18751
rect 7331 18717 7340 18751
rect 7288 18708 7340 18717
rect 7472 18708 7524 18760
rect 8208 18776 8260 18828
rect 3884 18640 3936 18692
rect 4344 18683 4396 18692
rect 4344 18649 4353 18683
rect 4353 18649 4387 18683
rect 4387 18649 4396 18683
rect 4344 18640 4396 18649
rect 4436 18683 4488 18692
rect 4436 18649 4445 18683
rect 4445 18649 4479 18683
rect 4479 18649 4488 18683
rect 4436 18640 4488 18649
rect 4620 18640 4672 18692
rect 6276 18640 6328 18692
rect 6736 18640 6788 18692
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 8944 18751 8996 18760
rect 8944 18717 8953 18751
rect 8953 18717 8987 18751
rect 8987 18717 8996 18751
rect 8944 18708 8996 18717
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 9128 18640 9180 18692
rect 9680 18640 9732 18692
rect 10140 18640 10192 18692
rect 10416 18708 10468 18760
rect 14372 18844 14424 18896
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14556 18708 14608 18760
rect 14740 18751 14792 18760
rect 14740 18717 14749 18751
rect 14749 18717 14783 18751
rect 14783 18717 14792 18751
rect 14740 18708 14792 18717
rect 17132 18844 17184 18896
rect 17776 18776 17828 18828
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 17132 18708 17184 18760
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 17408 18751 17460 18760
rect 17408 18717 17417 18751
rect 17417 18717 17451 18751
rect 17451 18717 17460 18751
rect 17408 18708 17460 18717
rect 17500 18708 17552 18760
rect 17684 18708 17736 18760
rect 17960 18751 18012 18760
rect 17960 18717 17969 18751
rect 17969 18717 18003 18751
rect 18003 18717 18012 18751
rect 17960 18708 18012 18717
rect 18880 18844 18932 18896
rect 20352 18844 20404 18896
rect 20076 18776 20128 18828
rect 21640 18776 21692 18828
rect 18972 18708 19024 18760
rect 19340 18708 19392 18760
rect 19984 18708 20036 18760
rect 21364 18751 21416 18760
rect 21364 18717 21373 18751
rect 21373 18717 21407 18751
rect 21407 18717 21416 18751
rect 21364 18708 21416 18717
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 22836 18751 22888 18760
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 27804 18751 27856 18760
rect 27804 18717 27813 18751
rect 27813 18717 27847 18751
rect 27847 18717 27856 18751
rect 27804 18708 27856 18717
rect 29092 18819 29144 18828
rect 29092 18785 29101 18819
rect 29101 18785 29135 18819
rect 29135 18785 29144 18819
rect 29092 18776 29144 18785
rect 29368 18751 29420 18760
rect 29368 18717 29377 18751
rect 29377 18717 29411 18751
rect 29411 18717 29420 18751
rect 29368 18708 29420 18717
rect 8300 18572 8352 18624
rect 10324 18572 10376 18624
rect 14924 18615 14976 18624
rect 14924 18581 14933 18615
rect 14933 18581 14967 18615
rect 14967 18581 14976 18615
rect 14924 18572 14976 18581
rect 15292 18683 15344 18692
rect 15292 18649 15301 18683
rect 15301 18649 15335 18683
rect 15335 18649 15344 18683
rect 15292 18640 15344 18649
rect 16764 18572 16816 18624
rect 16856 18615 16908 18624
rect 16856 18581 16865 18615
rect 16865 18581 16899 18615
rect 16899 18581 16908 18615
rect 16856 18572 16908 18581
rect 17040 18572 17092 18624
rect 18328 18683 18380 18692
rect 18328 18649 18337 18683
rect 18337 18649 18371 18683
rect 18371 18649 18380 18683
rect 18328 18640 18380 18649
rect 18880 18640 18932 18692
rect 26792 18640 26844 18692
rect 27160 18640 27212 18692
rect 27528 18683 27580 18692
rect 27528 18649 27537 18683
rect 27537 18649 27571 18683
rect 27571 18649 27580 18683
rect 27528 18640 27580 18649
rect 27896 18572 27948 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 2596 18368 2648 18420
rect 4436 18368 4488 18420
rect 10416 18300 10468 18352
rect 11060 18368 11112 18420
rect 12072 18368 12124 18420
rect 15292 18368 15344 18420
rect 17500 18411 17552 18420
rect 17500 18377 17509 18411
rect 17509 18377 17543 18411
rect 17543 18377 17552 18411
rect 17500 18368 17552 18377
rect 18328 18368 18380 18420
rect 18604 18368 18656 18420
rect 20076 18368 20128 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 21364 18368 21416 18420
rect 15200 18343 15252 18352
rect 15200 18309 15218 18343
rect 15218 18309 15252 18343
rect 1860 18232 1912 18284
rect 2136 18275 2188 18284
rect 2136 18241 2145 18275
rect 2145 18241 2179 18275
rect 2179 18241 2188 18275
rect 2136 18232 2188 18241
rect 3148 18232 3200 18284
rect 3332 18164 3384 18216
rect 4160 18232 4212 18284
rect 4620 18232 4672 18284
rect 5264 18232 5316 18284
rect 5448 18232 5500 18284
rect 15200 18300 15252 18309
rect 10968 18275 11020 18284
rect 10968 18241 10977 18275
rect 10977 18241 11011 18275
rect 11011 18241 11020 18275
rect 10968 18232 11020 18241
rect 11796 18275 11848 18284
rect 11796 18241 11805 18275
rect 11805 18241 11839 18275
rect 11839 18241 11848 18275
rect 11796 18232 11848 18241
rect 14280 18232 14332 18284
rect 5724 18164 5776 18216
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 10876 18164 10928 18216
rect 12072 18207 12124 18216
rect 12072 18173 12081 18207
rect 12081 18173 12115 18207
rect 12115 18173 12124 18207
rect 12072 18164 12124 18173
rect 16856 18300 16908 18352
rect 4252 18139 4304 18148
rect 4252 18105 4261 18139
rect 4261 18105 4295 18139
rect 4295 18105 4304 18139
rect 4252 18096 4304 18105
rect 5356 18096 5408 18148
rect 5540 18096 5592 18148
rect 8944 18096 8996 18148
rect 14924 18096 14976 18148
rect 15844 18232 15896 18284
rect 16764 18275 16816 18284
rect 16764 18241 16774 18275
rect 16774 18241 16808 18275
rect 16808 18241 16816 18275
rect 16764 18232 16816 18241
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17684 18275 17736 18284
rect 17684 18241 17693 18275
rect 17693 18241 17727 18275
rect 17727 18241 17736 18275
rect 17684 18232 17736 18241
rect 17960 18232 18012 18284
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 18420 18275 18472 18284
rect 18420 18241 18429 18275
rect 18429 18241 18463 18275
rect 18463 18241 18472 18275
rect 18420 18232 18472 18241
rect 10416 18028 10468 18080
rect 10784 18028 10836 18080
rect 12624 18028 12676 18080
rect 15660 18028 15712 18080
rect 16856 18096 16908 18148
rect 17684 18096 17736 18148
rect 17316 18071 17368 18080
rect 17316 18037 17325 18071
rect 17325 18037 17359 18071
rect 17359 18037 17368 18071
rect 17316 18028 17368 18037
rect 18512 18028 18564 18080
rect 18972 18232 19024 18284
rect 21180 18232 21232 18284
rect 21272 18232 21324 18284
rect 21548 18232 21600 18284
rect 21916 18275 21968 18284
rect 21916 18241 21925 18275
rect 21925 18241 21959 18275
rect 21959 18241 21968 18275
rect 21916 18232 21968 18241
rect 27528 18368 27580 18420
rect 24584 18300 24636 18352
rect 27896 18343 27948 18352
rect 27896 18309 27905 18343
rect 27905 18309 27939 18343
rect 27939 18309 27948 18343
rect 27896 18300 27948 18309
rect 28908 18300 28960 18352
rect 21640 18139 21692 18148
rect 21640 18105 21649 18139
rect 21649 18105 21683 18139
rect 21683 18105 21692 18139
rect 21640 18096 21692 18105
rect 22192 18096 22244 18148
rect 18788 18028 18840 18080
rect 22008 18028 22060 18080
rect 23296 18275 23348 18284
rect 23296 18241 23305 18275
rect 23305 18241 23339 18275
rect 23339 18241 23348 18275
rect 23296 18232 23348 18241
rect 25044 18164 25096 18216
rect 26240 18275 26292 18284
rect 26240 18241 26249 18275
rect 26249 18241 26283 18275
rect 26283 18241 26292 18275
rect 26240 18232 26292 18241
rect 27620 18275 27672 18284
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 26332 18164 26384 18216
rect 25504 18028 25556 18080
rect 26240 18028 26292 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2136 17824 2188 17876
rect 2504 17824 2556 17876
rect 3424 17824 3476 17876
rect 4068 17824 4120 17876
rect 4160 17756 4212 17808
rect 4344 17688 4396 17740
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 3148 17595 3200 17604
rect 3148 17561 3157 17595
rect 3157 17561 3191 17595
rect 3191 17561 3200 17595
rect 3148 17552 3200 17561
rect 3332 17663 3384 17672
rect 3332 17629 3341 17663
rect 3341 17629 3375 17663
rect 3375 17629 3384 17663
rect 3332 17620 3384 17629
rect 3424 17552 3476 17604
rect 3792 17620 3844 17672
rect 4160 17663 4212 17672
rect 4160 17629 4169 17663
rect 4169 17629 4203 17663
rect 4203 17629 4212 17663
rect 4160 17620 4212 17629
rect 4252 17663 4304 17672
rect 4252 17629 4261 17663
rect 4261 17629 4295 17663
rect 4295 17629 4304 17663
rect 4252 17620 4304 17629
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 5356 17756 5408 17808
rect 5724 17731 5776 17740
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 3884 17484 3936 17536
rect 4252 17484 4304 17536
rect 6276 17824 6328 17876
rect 8300 17824 8352 17876
rect 8944 17824 8996 17876
rect 10692 17824 10744 17876
rect 12072 17824 12124 17876
rect 18328 17824 18380 17876
rect 21916 17824 21968 17876
rect 24584 17824 24636 17876
rect 28908 17824 28960 17876
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 7564 17620 7616 17672
rect 8484 17620 8536 17672
rect 11060 17688 11112 17740
rect 6920 17552 6972 17604
rect 7840 17552 7892 17604
rect 7104 17484 7156 17536
rect 8392 17484 8444 17536
rect 9864 17552 9916 17604
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 10968 17620 11020 17672
rect 12532 17756 12584 17808
rect 13728 17756 13780 17808
rect 17960 17756 18012 17808
rect 18696 17756 18748 17808
rect 27436 17799 27488 17808
rect 27436 17765 27445 17799
rect 27445 17765 27479 17799
rect 27479 17765 27488 17799
rect 27436 17756 27488 17765
rect 11980 17688 12032 17740
rect 9128 17527 9180 17536
rect 9128 17493 9137 17527
rect 9137 17493 9171 17527
rect 9171 17493 9180 17527
rect 9128 17484 9180 17493
rect 10784 17484 10836 17536
rect 12072 17552 12124 17604
rect 12256 17552 12308 17604
rect 17316 17688 17368 17740
rect 19432 17688 19484 17740
rect 20260 17688 20312 17740
rect 22100 17688 22152 17740
rect 27620 17688 27672 17740
rect 15660 17663 15712 17672
rect 15660 17629 15669 17663
rect 15669 17629 15703 17663
rect 15703 17629 15712 17663
rect 15660 17620 15712 17629
rect 18420 17620 18472 17672
rect 21640 17620 21692 17672
rect 21824 17663 21876 17672
rect 21824 17629 21833 17663
rect 21833 17629 21867 17663
rect 21867 17629 21876 17663
rect 21824 17620 21876 17629
rect 12808 17552 12860 17604
rect 19984 17552 20036 17604
rect 11704 17484 11756 17536
rect 12348 17484 12400 17536
rect 15108 17484 15160 17536
rect 15292 17484 15344 17536
rect 19708 17484 19760 17536
rect 21272 17484 21324 17536
rect 24676 17620 24728 17672
rect 27528 17620 27580 17672
rect 25504 17595 25556 17604
rect 25504 17561 25513 17595
rect 25513 17561 25547 17595
rect 25547 17561 25556 17595
rect 25504 17552 25556 17561
rect 26240 17552 26292 17604
rect 26792 17552 26844 17604
rect 22100 17484 22152 17536
rect 26332 17484 26384 17536
rect 27160 17484 27212 17536
rect 27712 17484 27764 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 3332 17280 3384 17332
rect 848 17212 900 17264
rect 3700 17212 3752 17264
rect 4528 17280 4580 17332
rect 5724 17280 5776 17332
rect 6920 17323 6972 17332
rect 6920 17289 6929 17323
rect 6929 17289 6963 17323
rect 6963 17289 6972 17323
rect 6920 17280 6972 17289
rect 7104 17323 7156 17332
rect 7104 17289 7113 17323
rect 7113 17289 7147 17323
rect 7147 17289 7156 17323
rect 7104 17280 7156 17289
rect 7564 17280 7616 17332
rect 7656 17280 7708 17332
rect 10232 17280 10284 17332
rect 10416 17280 10468 17332
rect 10968 17280 11020 17332
rect 19708 17323 19760 17332
rect 19708 17289 19717 17323
rect 19717 17289 19751 17323
rect 19751 17289 19760 17323
rect 19708 17280 19760 17289
rect 19984 17280 20036 17332
rect 21364 17280 21416 17332
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 4344 17144 4396 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 8300 17187 8352 17196
rect 8300 17153 8309 17187
rect 8309 17153 8343 17187
rect 8343 17153 8352 17187
rect 8300 17144 8352 17153
rect 4712 17076 4764 17128
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 8392 17119 8444 17128
rect 8392 17085 8401 17119
rect 8401 17085 8435 17119
rect 8435 17085 8444 17119
rect 8392 17076 8444 17085
rect 4620 17008 4672 17060
rect 7840 17008 7892 17060
rect 9680 17144 9732 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 10600 17144 10652 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10968 17187 11020 17196
rect 10968 17153 10977 17187
rect 10977 17153 11011 17187
rect 11011 17153 11020 17187
rect 10968 17144 11020 17153
rect 11336 17187 11388 17196
rect 11336 17153 11345 17187
rect 11345 17153 11379 17187
rect 11379 17153 11388 17187
rect 11336 17144 11388 17153
rect 12808 17187 12860 17196
rect 12808 17153 12817 17187
rect 12817 17153 12851 17187
rect 12851 17153 12860 17187
rect 12808 17144 12860 17153
rect 13728 17144 13780 17196
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 14280 17076 14332 17128
rect 15016 17076 15068 17128
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 18420 17212 18472 17264
rect 19248 17212 19300 17264
rect 21548 17280 21600 17332
rect 21732 17212 21784 17264
rect 21364 17144 21416 17196
rect 21640 17187 21692 17196
rect 21640 17153 21649 17187
rect 21649 17153 21683 17187
rect 21683 17153 21692 17187
rect 21640 17144 21692 17153
rect 22100 17280 22152 17332
rect 27068 17280 27120 17332
rect 18144 17119 18196 17128
rect 18144 17085 18153 17119
rect 18153 17085 18187 17119
rect 18187 17085 18196 17119
rect 18144 17076 18196 17085
rect 12900 17008 12952 17060
rect 19432 17076 19484 17128
rect 21916 17187 21968 17196
rect 21916 17153 21926 17187
rect 21926 17153 21960 17187
rect 21960 17153 21968 17187
rect 21916 17144 21968 17153
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 26792 17255 26844 17264
rect 26792 17221 26801 17255
rect 26801 17221 26835 17255
rect 26835 17221 26844 17255
rect 26792 17212 26844 17221
rect 19800 17008 19852 17060
rect 12348 16940 12400 16992
rect 12716 16940 12768 16992
rect 16580 16940 16632 16992
rect 21640 16940 21692 16992
rect 25596 17187 25648 17196
rect 25596 17153 25605 17187
rect 25605 17153 25639 17187
rect 25639 17153 25648 17187
rect 25596 17144 25648 17153
rect 26332 17144 26384 17196
rect 27620 17212 27672 17264
rect 27712 17255 27764 17264
rect 27712 17221 27721 17255
rect 27721 17221 27755 17255
rect 27755 17221 27764 17255
rect 27712 17212 27764 17221
rect 28724 17212 28776 17264
rect 26056 17076 26108 17128
rect 22376 16940 22428 16992
rect 25412 16983 25464 16992
rect 25412 16949 25421 16983
rect 25421 16949 25455 16983
rect 25455 16949 25464 16983
rect 25412 16940 25464 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 17960 16736 18012 16788
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 21272 16736 21324 16788
rect 5724 16668 5776 16720
rect 2872 16600 2924 16652
rect 848 16532 900 16584
rect 6828 16600 6880 16652
rect 8392 16668 8444 16720
rect 8852 16600 8904 16652
rect 7288 16532 7340 16584
rect 8208 16532 8260 16584
rect 9864 16532 9916 16584
rect 10324 16600 10376 16652
rect 14648 16668 14700 16720
rect 17408 16668 17460 16720
rect 18052 16668 18104 16720
rect 24492 16668 24544 16720
rect 13452 16600 13504 16652
rect 16672 16600 16724 16652
rect 1584 16464 1636 16516
rect 7012 16464 7064 16516
rect 10968 16532 11020 16584
rect 12716 16575 12768 16584
rect 12716 16541 12725 16575
rect 12725 16541 12759 16575
rect 12759 16541 12768 16575
rect 12716 16532 12768 16541
rect 12900 16575 12952 16584
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 13084 16575 13136 16584
rect 13084 16541 13093 16575
rect 13093 16541 13127 16575
rect 13127 16541 13136 16575
rect 13084 16532 13136 16541
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 16580 16532 16632 16584
rect 17408 16575 17460 16584
rect 17408 16541 17417 16575
rect 17417 16541 17451 16575
rect 17451 16541 17460 16575
rect 17408 16532 17460 16541
rect 6644 16439 6696 16448
rect 6644 16405 6653 16439
rect 6653 16405 6687 16439
rect 6687 16405 6696 16439
rect 6644 16396 6696 16405
rect 10048 16396 10100 16448
rect 13728 16464 13780 16516
rect 15476 16507 15528 16516
rect 15476 16473 15485 16507
rect 15485 16473 15519 16507
rect 15519 16473 15528 16507
rect 15476 16464 15528 16473
rect 17868 16532 17920 16584
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 17960 16532 18012 16541
rect 18052 16532 18104 16584
rect 20260 16600 20312 16652
rect 21180 16600 21232 16652
rect 21364 16600 21416 16652
rect 19708 16532 19760 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 21640 16575 21692 16584
rect 21640 16541 21649 16575
rect 21649 16541 21683 16575
rect 21683 16541 21692 16575
rect 21640 16532 21692 16541
rect 20352 16464 20404 16516
rect 21548 16464 21600 16516
rect 21824 16532 21876 16584
rect 22376 16643 22428 16652
rect 22376 16609 22385 16643
rect 22385 16609 22419 16643
rect 22419 16609 22428 16643
rect 22376 16600 22428 16609
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 24676 16532 24728 16584
rect 25596 16736 25648 16788
rect 27436 16736 27488 16788
rect 28724 16736 28776 16788
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 26056 16600 26108 16652
rect 27068 16643 27120 16652
rect 27068 16609 27077 16643
rect 27077 16609 27111 16643
rect 27111 16609 27120 16643
rect 27068 16600 27120 16609
rect 27160 16643 27212 16652
rect 27160 16609 27169 16643
rect 27169 16609 27203 16643
rect 27203 16609 27212 16643
rect 27160 16600 27212 16609
rect 29092 16711 29144 16720
rect 29092 16677 29101 16711
rect 29101 16677 29135 16711
rect 29135 16677 29144 16711
rect 29092 16668 29144 16677
rect 27436 16600 27488 16652
rect 28172 16532 28224 16584
rect 29276 16575 29328 16584
rect 29276 16541 29285 16575
rect 29285 16541 29319 16575
rect 29319 16541 29328 16575
rect 29276 16532 29328 16541
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 13544 16396 13596 16448
rect 14280 16396 14332 16448
rect 17500 16439 17552 16448
rect 17500 16405 17509 16439
rect 17509 16405 17543 16439
rect 17543 16405 17552 16439
rect 17500 16396 17552 16405
rect 17776 16396 17828 16448
rect 17868 16396 17920 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 22100 16396 22152 16448
rect 24032 16396 24084 16448
rect 25044 16439 25096 16448
rect 25044 16405 25053 16439
rect 25053 16405 25087 16439
rect 25087 16405 25096 16439
rect 25044 16396 25096 16405
rect 25504 16464 25556 16516
rect 26424 16464 26476 16516
rect 26056 16396 26108 16448
rect 28448 16439 28500 16448
rect 28448 16405 28457 16439
rect 28457 16405 28491 16439
rect 28491 16405 28500 16439
rect 28448 16396 28500 16405
rect 28908 16439 28960 16448
rect 28908 16405 28917 16439
rect 28917 16405 28951 16439
rect 28951 16405 28960 16439
rect 28908 16396 28960 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 6000 16192 6052 16244
rect 2596 16124 2648 16176
rect 3792 16124 3844 16176
rect 3332 16056 3384 16108
rect 3884 16056 3936 16108
rect 4712 16124 4764 16176
rect 5448 16124 5500 16176
rect 9128 16192 9180 16244
rect 10324 16192 10376 16244
rect 11704 16192 11756 16244
rect 12072 16192 12124 16244
rect 13728 16192 13780 16244
rect 6644 16124 6696 16176
rect 8208 16124 8260 16176
rect 9036 16124 9088 16176
rect 4252 16056 4304 16108
rect 3608 15988 3660 16040
rect 4620 16099 4672 16108
rect 4620 16065 4629 16099
rect 4629 16065 4663 16099
rect 4663 16065 4672 16099
rect 4620 16056 4672 16065
rect 3976 15920 4028 15972
rect 5172 16099 5224 16108
rect 5172 16065 5181 16099
rect 5181 16065 5215 16099
rect 5215 16065 5224 16099
rect 5172 16056 5224 16065
rect 5356 16099 5408 16108
rect 5356 16065 5365 16099
rect 5365 16065 5399 16099
rect 5399 16065 5408 16099
rect 5356 16056 5408 16065
rect 6000 16056 6052 16108
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 5632 15988 5684 16040
rect 6644 16031 6696 16040
rect 6644 15997 6653 16031
rect 6653 15997 6687 16031
rect 6687 15997 6696 16031
rect 6644 15988 6696 15997
rect 8944 16031 8996 16040
rect 8944 15997 8953 16031
rect 8953 15997 8987 16031
rect 8987 15997 8996 16031
rect 8944 15988 8996 15997
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 10048 16099 10100 16108
rect 10048 16065 10057 16099
rect 10057 16065 10091 16099
rect 10091 16065 10100 16099
rect 10048 16056 10100 16065
rect 5724 15920 5776 15972
rect 10048 15920 10100 15972
rect 4620 15852 4672 15904
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 9864 15852 9916 15904
rect 10324 15920 10376 15972
rect 10784 16056 10836 16108
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11796 16124 11848 16176
rect 13452 16124 13504 16176
rect 13544 16167 13596 16176
rect 13544 16133 13553 16167
rect 13553 16133 13587 16167
rect 13587 16133 13596 16167
rect 13544 16124 13596 16133
rect 14280 16124 14332 16176
rect 15476 16192 15528 16244
rect 16672 16192 16724 16244
rect 18696 16192 18748 16244
rect 19616 16192 19668 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 17776 16124 17828 16176
rect 10508 15988 10560 16040
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 19340 16056 19392 16108
rect 19708 16099 19760 16108
rect 19708 16065 19717 16099
rect 19717 16065 19751 16099
rect 19751 16065 19760 16099
rect 19708 16056 19760 16065
rect 14280 15988 14332 16040
rect 16120 16031 16172 16040
rect 16120 15997 16129 16031
rect 16129 15997 16163 16031
rect 16163 15997 16172 16031
rect 16120 15988 16172 15997
rect 17592 15988 17644 16040
rect 17868 15988 17920 16040
rect 18144 15988 18196 16040
rect 19248 15988 19300 16040
rect 12900 15920 12952 15972
rect 17500 15920 17552 15972
rect 17960 15920 18012 15972
rect 18880 15920 18932 15972
rect 19432 15988 19484 16040
rect 20260 16099 20312 16108
rect 20260 16065 20291 16099
rect 20291 16065 20312 16099
rect 20260 16056 20312 16065
rect 20352 16099 20404 16108
rect 20352 16065 20361 16099
rect 20361 16065 20395 16099
rect 20395 16065 20404 16099
rect 20352 16056 20404 16065
rect 20904 16056 20956 16108
rect 22468 16192 22520 16244
rect 24676 16192 24728 16244
rect 25504 16192 25556 16244
rect 26424 16192 26476 16244
rect 24032 16124 24084 16176
rect 24492 16167 24544 16176
rect 24492 16133 24501 16167
rect 24501 16133 24535 16167
rect 24535 16133 24544 16167
rect 24492 16124 24544 16133
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 25044 16056 25096 16108
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 27436 16124 27488 16176
rect 26240 16056 26292 16108
rect 27896 16192 27948 16244
rect 28908 16124 28960 16176
rect 21180 15988 21232 16040
rect 22008 15988 22060 16040
rect 25136 15988 25188 16040
rect 27252 16031 27304 16040
rect 27252 15997 27261 16031
rect 27261 15997 27295 16031
rect 27295 15997 27304 16031
rect 27252 15988 27304 15997
rect 27620 16031 27672 16040
rect 27620 15997 27629 16031
rect 27629 15997 27663 16031
rect 27663 15997 27672 16031
rect 27620 15988 27672 15997
rect 20260 15920 20312 15972
rect 21916 15920 21968 15972
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 15660 15852 15712 15904
rect 16396 15852 16448 15904
rect 19432 15852 19484 15904
rect 19616 15852 19668 15904
rect 22100 15895 22152 15904
rect 22100 15861 22109 15895
rect 22109 15861 22143 15895
rect 22143 15861 22152 15895
rect 22100 15852 22152 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2596 15691 2648 15700
rect 2596 15657 2605 15691
rect 2605 15657 2639 15691
rect 2639 15657 2648 15691
rect 2596 15648 2648 15657
rect 3608 15691 3660 15700
rect 3608 15657 3617 15691
rect 3617 15657 3651 15691
rect 3651 15657 3660 15691
rect 3608 15648 3660 15657
rect 3700 15648 3752 15700
rect 4068 15648 4120 15700
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2872 15444 2924 15496
rect 3332 15444 3384 15496
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4068 15444 4120 15496
rect 4620 15444 4672 15496
rect 5172 15512 5224 15564
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 6644 15648 6696 15700
rect 8944 15648 8996 15700
rect 10048 15648 10100 15700
rect 10324 15648 10376 15700
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 10968 15648 11020 15700
rect 11796 15691 11848 15700
rect 11796 15657 11805 15691
rect 11805 15657 11839 15691
rect 11839 15657 11848 15691
rect 11796 15648 11848 15657
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 16488 15648 16540 15700
rect 18236 15648 18288 15700
rect 12072 15580 12124 15632
rect 7656 15512 7708 15564
rect 9772 15512 9824 15564
rect 12900 15512 12952 15564
rect 1492 15419 1544 15428
rect 1492 15385 1501 15419
rect 1501 15385 1535 15419
rect 1535 15385 1544 15419
rect 1492 15376 1544 15385
rect 8484 15444 8536 15496
rect 9036 15444 9088 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 10232 15444 10284 15496
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11336 15444 11388 15496
rect 12992 15487 13044 15496
rect 12992 15453 13001 15487
rect 13001 15453 13035 15487
rect 13035 15453 13044 15487
rect 12992 15444 13044 15453
rect 13176 15444 13228 15496
rect 14004 15512 14056 15564
rect 5632 15376 5684 15428
rect 7288 15376 7340 15428
rect 9864 15376 9916 15428
rect 14372 15444 14424 15496
rect 15292 15512 15344 15564
rect 15660 15512 15712 15564
rect 17776 15512 17828 15564
rect 17960 15555 18012 15564
rect 17960 15521 17969 15555
rect 17969 15521 18003 15555
rect 18003 15521 18012 15555
rect 17960 15512 18012 15521
rect 18880 15648 18932 15700
rect 20352 15648 20404 15700
rect 21272 15648 21324 15700
rect 19892 15512 19944 15564
rect 22284 15580 22336 15632
rect 23572 15512 23624 15564
rect 16304 15444 16356 15496
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 9772 15308 9824 15360
rect 12624 15351 12676 15360
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 13084 15308 13136 15360
rect 14280 15308 14332 15360
rect 15292 15376 15344 15428
rect 18236 15376 18288 15428
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 19524 15444 19576 15496
rect 20720 15487 20772 15496
rect 20720 15453 20729 15487
rect 20729 15453 20763 15487
rect 20763 15453 20772 15487
rect 20720 15444 20772 15453
rect 22376 15444 22428 15496
rect 23664 15487 23716 15496
rect 22008 15376 22060 15428
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 24676 15444 24728 15496
rect 27344 15487 27396 15496
rect 27344 15453 27353 15487
rect 27353 15453 27387 15487
rect 27387 15453 27396 15487
rect 27344 15444 27396 15453
rect 22468 15308 22520 15360
rect 27160 15376 27212 15428
rect 29092 15487 29144 15496
rect 29092 15453 29101 15487
rect 29101 15453 29135 15487
rect 29135 15453 29144 15487
rect 29092 15444 29144 15453
rect 29368 15487 29420 15496
rect 29368 15453 29377 15487
rect 29377 15453 29411 15487
rect 29411 15453 29420 15487
rect 29368 15444 29420 15453
rect 23204 15351 23256 15360
rect 23204 15317 23213 15351
rect 23213 15317 23247 15351
rect 23247 15317 23256 15351
rect 23204 15308 23256 15317
rect 24400 15308 24452 15360
rect 27252 15308 27304 15360
rect 28540 15308 28592 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 4068 15104 4120 15156
rect 9680 15104 9732 15156
rect 10140 15104 10192 15156
rect 11612 15104 11664 15156
rect 12348 15104 12400 15156
rect 12624 15104 12676 15156
rect 12992 15104 13044 15156
rect 17316 15104 17368 15156
rect 19248 15104 19300 15156
rect 20904 15104 20956 15156
rect 23664 15104 23716 15156
rect 27896 15147 27948 15156
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 7840 15036 7892 15088
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 11152 14968 11204 15020
rect 11612 14968 11664 15020
rect 12348 15011 12400 15020
rect 12348 14977 12357 15011
rect 12357 14977 12391 15011
rect 12391 14977 12400 15011
rect 12348 14968 12400 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 8300 14900 8352 14952
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 16212 15036 16264 15088
rect 16304 15079 16356 15088
rect 16304 15045 16313 15079
rect 16313 15045 16347 15079
rect 16347 15045 16356 15079
rect 16304 15036 16356 15045
rect 19340 15036 19392 15088
rect 23204 15036 23256 15088
rect 1952 14832 2004 14884
rect 9128 14832 9180 14884
rect 11888 14875 11940 14884
rect 11888 14841 11897 14875
rect 11897 14841 11931 14875
rect 11931 14841 11940 14875
rect 11888 14832 11940 14841
rect 13084 14900 13136 14952
rect 14280 14943 14332 14952
rect 14280 14909 14289 14943
rect 14289 14909 14323 14943
rect 14323 14909 14332 14943
rect 14280 14900 14332 14909
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 17408 14968 17460 15020
rect 22008 15011 22060 15020
rect 22008 14977 22017 15011
rect 22017 14977 22051 15011
rect 22051 14977 22060 15011
rect 22008 14968 22060 14977
rect 24400 14968 24452 15020
rect 26240 14968 26292 15020
rect 27896 15113 27905 15147
rect 27905 15113 27939 15147
rect 27939 15113 27948 15147
rect 27896 15104 27948 15113
rect 27988 15104 28040 15156
rect 20904 14900 20956 14952
rect 22284 14900 22336 14952
rect 25136 14900 25188 14952
rect 26056 14900 26108 14952
rect 12440 14832 12492 14884
rect 13544 14832 13596 14884
rect 14096 14832 14148 14884
rect 6736 14807 6788 14816
rect 6736 14773 6745 14807
rect 6745 14773 6779 14807
rect 6779 14773 6788 14807
rect 6736 14764 6788 14773
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 10140 14764 10192 14816
rect 13268 14764 13320 14816
rect 13360 14764 13412 14816
rect 22928 14832 22980 14884
rect 18236 14764 18288 14816
rect 20444 14764 20496 14816
rect 22100 14764 22152 14816
rect 25412 14807 25464 14816
rect 25412 14773 25421 14807
rect 25421 14773 25455 14807
rect 25455 14773 25464 14807
rect 25412 14764 25464 14773
rect 26240 14764 26292 14816
rect 27160 14943 27212 14952
rect 27160 14909 27169 14943
rect 27169 14909 27203 14943
rect 27203 14909 27212 14943
rect 27160 14900 27212 14909
rect 27344 14943 27396 14952
rect 27344 14909 27353 14943
rect 27353 14909 27387 14943
rect 27387 14909 27396 14943
rect 27344 14900 27396 14909
rect 27436 14943 27488 14952
rect 27436 14909 27445 14943
rect 27445 14909 27479 14943
rect 27479 14909 27488 14943
rect 27436 14900 27488 14909
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 28172 14875 28224 14884
rect 28172 14841 28181 14875
rect 28181 14841 28215 14875
rect 28215 14841 28224 14875
rect 28172 14832 28224 14841
rect 28264 14807 28316 14816
rect 28264 14773 28273 14807
rect 28273 14773 28307 14807
rect 28307 14773 28316 14807
rect 28264 14764 28316 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 6736 14603 6788 14612
rect 6736 14569 6745 14603
rect 6745 14569 6779 14603
rect 6779 14569 6788 14603
rect 6736 14560 6788 14569
rect 6828 14560 6880 14612
rect 6920 14492 6972 14544
rect 4804 14424 4856 14476
rect 7380 14424 7432 14476
rect 8484 14424 8536 14476
rect 2780 14356 2832 14408
rect 6000 14356 6052 14408
rect 6828 14356 6880 14408
rect 14188 14560 14240 14612
rect 14556 14560 14608 14612
rect 15936 14603 15988 14612
rect 15936 14569 15945 14603
rect 15945 14569 15979 14603
rect 15979 14569 15988 14603
rect 15936 14560 15988 14569
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 10048 14492 10100 14544
rect 10324 14492 10376 14544
rect 10600 14492 10652 14544
rect 9220 14424 9272 14476
rect 10784 14424 10836 14476
rect 11244 14492 11296 14544
rect 17960 14535 18012 14544
rect 17960 14501 17969 14535
rect 17969 14501 18003 14535
rect 18003 14501 18012 14535
rect 17960 14492 18012 14501
rect 18236 14492 18288 14544
rect 18512 14492 18564 14544
rect 19524 14492 19576 14544
rect 10048 14399 10100 14408
rect 10048 14365 10057 14399
rect 10057 14365 10091 14399
rect 10091 14365 10100 14399
rect 10048 14356 10100 14365
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 10600 14399 10652 14408
rect 10600 14365 10609 14399
rect 10609 14365 10643 14399
rect 10643 14365 10652 14399
rect 10600 14356 10652 14365
rect 11060 14356 11112 14408
rect 13084 14356 13136 14408
rect 14004 14424 14056 14476
rect 14188 14424 14240 14476
rect 15016 14424 15068 14476
rect 16396 14424 16448 14476
rect 4712 14331 4764 14340
rect 4712 14297 4721 14331
rect 4721 14297 4755 14331
rect 4755 14297 4764 14331
rect 4712 14288 4764 14297
rect 5448 14288 5500 14340
rect 3424 14220 3476 14272
rect 5540 14220 5592 14272
rect 6368 14288 6420 14340
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 11520 14288 11572 14340
rect 12992 14288 13044 14340
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 14372 14356 14424 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 15200 14356 15252 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 18604 14467 18656 14476
rect 18604 14433 18613 14467
rect 18613 14433 18647 14467
rect 18647 14433 18656 14467
rect 18604 14424 18656 14433
rect 20076 14424 20128 14476
rect 25136 14424 25188 14476
rect 27436 14560 27488 14612
rect 27712 14560 27764 14612
rect 28264 14560 28316 14612
rect 29092 14424 29144 14476
rect 14556 14288 14608 14340
rect 15016 14288 15068 14340
rect 17040 14288 17092 14340
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 10600 14220 10652 14272
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 13636 14220 13688 14272
rect 17408 14220 17460 14272
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 18512 14356 18564 14408
rect 18880 14356 18932 14408
rect 18328 14288 18380 14340
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 26240 14356 26292 14408
rect 27620 14399 27672 14408
rect 27620 14365 27629 14399
rect 27629 14365 27663 14399
rect 27663 14365 27672 14399
rect 27620 14356 27672 14365
rect 19984 14331 20036 14340
rect 19984 14297 19993 14331
rect 19993 14297 20027 14331
rect 20027 14297 20036 14331
rect 19984 14288 20036 14297
rect 20996 14288 21048 14340
rect 18236 14220 18288 14272
rect 20260 14220 20312 14272
rect 25412 14288 25464 14340
rect 27160 14331 27212 14340
rect 27160 14297 27169 14331
rect 27169 14297 27203 14331
rect 27203 14297 27212 14331
rect 27160 14288 27212 14297
rect 27344 14331 27396 14340
rect 27344 14297 27353 14331
rect 27353 14297 27387 14331
rect 27387 14297 27396 14331
rect 27344 14288 27396 14297
rect 28172 14288 28224 14340
rect 28908 14288 28960 14340
rect 22284 14220 22336 14272
rect 29184 14220 29236 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 1952 13812 2004 13864
rect 4804 14016 4856 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 6184 14016 6236 14068
rect 3424 13948 3476 14000
rect 5540 13948 5592 14000
rect 7012 14016 7064 14068
rect 10324 14016 10376 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 6920 13948 6972 14000
rect 4620 13880 4672 13932
rect 5448 13880 5500 13932
rect 6000 13880 6052 13932
rect 6828 13923 6880 13932
rect 6828 13889 6837 13923
rect 6837 13889 6871 13923
rect 6871 13889 6880 13923
rect 6828 13880 6880 13889
rect 4068 13812 4120 13864
rect 4712 13812 4764 13864
rect 7196 13812 7248 13864
rect 8300 13880 8352 13932
rect 9128 13923 9180 13932
rect 9128 13889 9137 13923
rect 9137 13889 9171 13923
rect 9171 13889 9180 13923
rect 9128 13880 9180 13889
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 3792 13676 3844 13728
rect 4068 13676 4120 13728
rect 7104 13676 7156 13728
rect 8208 13744 8260 13796
rect 11244 13948 11296 14000
rect 10508 13880 10560 13932
rect 10784 13923 10836 13932
rect 10784 13889 10791 13923
rect 10791 13889 10836 13923
rect 10784 13880 10836 13889
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11060 13880 11112 13932
rect 11612 13948 11664 14000
rect 13084 13991 13136 14000
rect 13084 13957 13093 13991
rect 13093 13957 13127 13991
rect 13127 13957 13136 13991
rect 13084 13948 13136 13957
rect 11520 13923 11572 13932
rect 11520 13889 11529 13923
rect 11529 13889 11563 13923
rect 11563 13889 11572 13923
rect 11520 13880 11572 13889
rect 10416 13744 10468 13796
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 12440 13812 12492 13864
rect 12992 13880 13044 13932
rect 13360 13923 13412 13932
rect 10968 13744 11020 13796
rect 13084 13812 13136 13864
rect 13360 13889 13368 13923
rect 13368 13889 13402 13923
rect 13402 13889 13412 13923
rect 13360 13880 13412 13889
rect 13636 13880 13688 13932
rect 13820 13948 13872 14000
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 14096 13880 14148 13932
rect 14556 13948 14608 14000
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 19432 14016 19484 14068
rect 19984 14016 20036 14068
rect 20076 14016 20128 14068
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 20996 14016 21048 14068
rect 22928 14016 22980 14068
rect 16028 13880 16080 13932
rect 17040 13880 17092 13932
rect 18144 13880 18196 13932
rect 18236 13923 18288 13932
rect 18236 13889 18245 13923
rect 18245 13889 18279 13923
rect 18279 13889 18288 13923
rect 18236 13880 18288 13889
rect 13544 13855 13596 13864
rect 13544 13821 13553 13855
rect 13553 13821 13587 13855
rect 13587 13821 13596 13855
rect 13544 13812 13596 13821
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 18696 13923 18748 13932
rect 18696 13889 18705 13923
rect 18705 13889 18739 13923
rect 18739 13889 18748 13923
rect 18696 13880 18748 13889
rect 19340 13812 19392 13864
rect 20628 13948 20680 14000
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 23480 13948 23532 14000
rect 28908 14059 28960 14068
rect 28908 14025 28917 14059
rect 28917 14025 28951 14059
rect 28951 14025 28960 14059
rect 28908 14016 28960 14025
rect 14648 13744 14700 13796
rect 19432 13744 19484 13796
rect 19800 13744 19852 13796
rect 19984 13744 20036 13796
rect 22008 13855 22060 13864
rect 22008 13821 22017 13855
rect 22017 13821 22051 13855
rect 22051 13821 22060 13855
rect 22008 13812 22060 13821
rect 26056 13880 26108 13932
rect 28816 13880 28868 13932
rect 29276 13923 29328 13932
rect 29276 13889 29285 13923
rect 29285 13889 29319 13923
rect 29319 13889 29328 13923
rect 29276 13880 29328 13889
rect 23204 13812 23256 13864
rect 9036 13719 9088 13728
rect 9036 13685 9045 13719
rect 9045 13685 9079 13719
rect 9079 13685 9088 13719
rect 9036 13676 9088 13685
rect 10508 13676 10560 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 11612 13676 11664 13728
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 12808 13719 12860 13728
rect 12808 13685 12817 13719
rect 12817 13685 12851 13719
rect 12851 13685 12860 13719
rect 12808 13676 12860 13685
rect 15660 13719 15712 13728
rect 15660 13685 15669 13719
rect 15669 13685 15703 13719
rect 15703 13685 15712 13719
rect 15660 13676 15712 13685
rect 16764 13719 16816 13728
rect 16764 13685 16773 13719
rect 16773 13685 16807 13719
rect 16807 13685 16816 13719
rect 16764 13676 16816 13685
rect 22284 13744 22336 13796
rect 22100 13676 22152 13728
rect 24952 13855 25004 13864
rect 24952 13821 24961 13855
rect 24961 13821 24995 13855
rect 24995 13821 25004 13855
rect 24952 13812 25004 13821
rect 27160 13855 27212 13864
rect 27160 13821 27169 13855
rect 27169 13821 27203 13855
rect 27203 13821 27212 13855
rect 27160 13812 27212 13821
rect 27528 13787 27580 13796
rect 27528 13753 27537 13787
rect 27537 13753 27571 13787
rect 27571 13753 27580 13787
rect 27528 13744 27580 13753
rect 25136 13676 25188 13728
rect 26424 13719 26476 13728
rect 26424 13685 26433 13719
rect 26433 13685 26467 13719
rect 26467 13685 26476 13719
rect 26424 13676 26476 13685
rect 27896 13676 27948 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 3792 13515 3844 13524
rect 3792 13481 3801 13515
rect 3801 13481 3835 13515
rect 3835 13481 3844 13515
rect 3792 13472 3844 13481
rect 11336 13472 11388 13524
rect 11796 13472 11848 13524
rect 19432 13472 19484 13524
rect 20444 13515 20496 13524
rect 20444 13481 20453 13515
rect 20453 13481 20487 13515
rect 20487 13481 20496 13515
rect 20444 13472 20496 13481
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 26056 13472 26108 13524
rect 27160 13472 27212 13524
rect 2596 13379 2648 13388
rect 2596 13345 2605 13379
rect 2605 13345 2639 13379
rect 2639 13345 2648 13379
rect 2596 13336 2648 13345
rect 4712 13336 4764 13388
rect 2504 13268 2556 13320
rect 3516 13268 3568 13320
rect 4068 13268 4120 13320
rect 7196 13268 7248 13320
rect 7656 13311 7708 13320
rect 7656 13277 7665 13311
rect 7665 13277 7699 13311
rect 7699 13277 7708 13311
rect 7656 13268 7708 13277
rect 7932 13311 7984 13320
rect 7932 13277 7941 13311
rect 7941 13277 7975 13311
rect 7975 13277 7984 13311
rect 7932 13268 7984 13277
rect 8116 13268 8168 13320
rect 11244 13336 11296 13388
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 2136 13175 2188 13184
rect 2136 13141 2145 13175
rect 2145 13141 2179 13175
rect 2179 13141 2188 13175
rect 2136 13132 2188 13141
rect 6276 13243 6328 13252
rect 6276 13209 6285 13243
rect 6285 13209 6319 13243
rect 6319 13209 6328 13243
rect 6276 13200 6328 13209
rect 6552 13200 6604 13252
rect 7288 13200 7340 13252
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 7564 13132 7616 13184
rect 7748 13132 7800 13184
rect 8484 13200 8536 13252
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 12072 13268 12124 13320
rect 12440 13404 12492 13456
rect 22008 13404 22060 13456
rect 14280 13336 14332 13388
rect 15660 13336 15712 13388
rect 16028 13336 16080 13388
rect 18236 13336 18288 13388
rect 18696 13336 18748 13388
rect 12808 13268 12860 13320
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 17132 13268 17184 13320
rect 11612 13243 11664 13252
rect 11612 13209 11621 13243
rect 11621 13209 11655 13243
rect 11655 13209 11664 13243
rect 11612 13200 11664 13209
rect 16764 13200 16816 13252
rect 19340 13268 19392 13320
rect 20444 13200 20496 13252
rect 9496 13132 9548 13184
rect 12900 13132 12952 13184
rect 17684 13132 17736 13184
rect 20628 13311 20680 13320
rect 20628 13277 20637 13311
rect 20637 13277 20671 13311
rect 20671 13277 20680 13311
rect 20628 13268 20680 13277
rect 25136 13336 25188 13388
rect 27620 13404 27672 13456
rect 27896 13379 27948 13388
rect 27896 13345 27905 13379
rect 27905 13345 27939 13379
rect 27939 13345 27948 13379
rect 27896 13336 27948 13345
rect 26332 13268 26384 13320
rect 26884 13268 26936 13320
rect 27160 13268 27212 13320
rect 20904 13243 20956 13252
rect 20904 13209 20913 13243
rect 20913 13209 20947 13243
rect 20947 13209 20956 13243
rect 20904 13200 20956 13209
rect 21916 13200 21968 13252
rect 24216 13200 24268 13252
rect 27068 13200 27120 13252
rect 27620 13311 27672 13320
rect 27620 13277 27629 13311
rect 27629 13277 27663 13311
rect 27663 13277 27672 13311
rect 27620 13268 27672 13277
rect 20720 13132 20772 13184
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 26608 13132 26660 13184
rect 27252 13132 27304 13184
rect 27712 13132 27764 13184
rect 28908 13200 28960 13252
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 3792 12928 3844 12980
rect 1952 12860 2004 12912
rect 2136 12860 2188 12912
rect 4068 12792 4120 12844
rect 4804 12860 4856 12912
rect 5540 12860 5592 12912
rect 6828 12928 6880 12980
rect 6276 12860 6328 12912
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 6736 12792 6788 12844
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7288 12792 7340 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 6000 12724 6052 12776
rect 7012 12724 7064 12776
rect 4620 12588 4672 12640
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 7840 12928 7892 12980
rect 7932 12928 7984 12980
rect 7932 12792 7984 12844
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 7656 12588 7708 12640
rect 7840 12588 7892 12640
rect 8208 12656 8260 12708
rect 10324 12928 10376 12980
rect 10232 12860 10284 12912
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 9036 12792 9088 12844
rect 8944 12724 8996 12776
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 11428 12792 11480 12844
rect 14280 12792 14332 12844
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 15844 12860 15896 12912
rect 17868 12928 17920 12980
rect 17684 12860 17736 12912
rect 19708 12928 19760 12980
rect 20628 12928 20680 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 24952 12928 25004 12980
rect 21272 12903 21324 12912
rect 21272 12869 21281 12903
rect 21281 12869 21315 12903
rect 21315 12869 21324 12903
rect 21272 12860 21324 12869
rect 22376 12860 22428 12912
rect 20444 12792 20496 12844
rect 20996 12792 21048 12844
rect 22008 12835 22060 12844
rect 22008 12801 22017 12835
rect 22017 12801 22051 12835
rect 22051 12801 22060 12835
rect 22008 12792 22060 12801
rect 26424 12928 26476 12980
rect 27160 12928 27212 12980
rect 27528 12971 27580 12980
rect 27528 12937 27537 12971
rect 27537 12937 27571 12971
rect 27571 12937 27580 12971
rect 27528 12928 27580 12937
rect 28908 12928 28960 12980
rect 26608 12835 26660 12844
rect 26608 12801 26617 12835
rect 26617 12801 26651 12835
rect 26651 12801 26660 12835
rect 26608 12792 26660 12801
rect 10416 12724 10468 12776
rect 10232 12656 10284 12708
rect 10784 12656 10836 12708
rect 11520 12656 11572 12708
rect 13084 12656 13136 12708
rect 13636 12656 13688 12708
rect 8944 12588 8996 12640
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 14924 12588 14976 12640
rect 16948 12767 17000 12776
rect 16948 12733 16957 12767
rect 16957 12733 16991 12767
rect 16991 12733 17000 12767
rect 16948 12724 17000 12733
rect 18880 12767 18932 12776
rect 18880 12733 18889 12767
rect 18889 12733 18923 12767
rect 18923 12733 18932 12767
rect 18880 12724 18932 12733
rect 22100 12724 22152 12776
rect 23664 12724 23716 12776
rect 27068 12835 27120 12844
rect 27068 12801 27077 12835
rect 27077 12801 27111 12835
rect 27111 12801 27120 12835
rect 27068 12792 27120 12801
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 27436 12792 27488 12844
rect 27988 12835 28040 12844
rect 27988 12801 27997 12835
rect 27997 12801 28031 12835
rect 28031 12801 28040 12835
rect 27988 12792 28040 12801
rect 28816 12792 28868 12844
rect 29276 12835 29328 12844
rect 29276 12801 29285 12835
rect 29285 12801 29319 12835
rect 29319 12801 29328 12835
rect 29276 12792 29328 12801
rect 27712 12724 27764 12776
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 25688 12631 25740 12640
rect 25688 12597 25697 12631
rect 25697 12597 25731 12631
rect 25731 12597 25740 12631
rect 25688 12588 25740 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 1676 12384 1728 12436
rect 2504 12384 2556 12436
rect 3332 12316 3384 12368
rect 4712 12316 4764 12368
rect 5540 12384 5592 12436
rect 6000 12427 6052 12436
rect 6000 12393 6009 12427
rect 6009 12393 6043 12427
rect 6043 12393 6052 12427
rect 6000 12384 6052 12393
rect 6644 12384 6696 12436
rect 7288 12384 7340 12436
rect 7472 12384 7524 12436
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 8760 12384 8812 12436
rect 10048 12427 10100 12436
rect 10048 12393 10057 12427
rect 10057 12393 10091 12427
rect 10091 12393 10100 12427
rect 10048 12384 10100 12393
rect 3976 12248 4028 12300
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 848 12180 900 12232
rect 3148 12180 3200 12232
rect 3424 12180 3476 12232
rect 5448 12316 5500 12368
rect 6552 12248 6604 12300
rect 10508 12427 10560 12436
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 11060 12384 11112 12436
rect 11244 12384 11296 12436
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 12532 12384 12584 12436
rect 6092 12180 6144 12232
rect 1952 12112 2004 12164
rect 6276 12180 6328 12232
rect 7932 12248 7984 12300
rect 9588 12248 9640 12300
rect 13268 12316 13320 12368
rect 14832 12384 14884 12436
rect 15844 12384 15896 12436
rect 16948 12384 17000 12436
rect 18880 12384 18932 12436
rect 27436 12384 27488 12436
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 7748 12180 7800 12232
rect 8116 12180 8168 12232
rect 8300 12180 8352 12232
rect 6368 12155 6420 12164
rect 6368 12121 6377 12155
rect 6377 12121 6411 12155
rect 6411 12121 6420 12155
rect 9680 12180 9732 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10232 12180 10284 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 6368 12112 6420 12121
rect 8944 12112 8996 12164
rect 10692 12155 10744 12164
rect 10692 12121 10701 12155
rect 10701 12121 10735 12155
rect 10735 12121 10744 12155
rect 10692 12112 10744 12121
rect 2228 12087 2280 12096
rect 2228 12053 2237 12087
rect 2237 12053 2271 12087
rect 2271 12053 2280 12087
rect 2228 12044 2280 12053
rect 7840 12044 7892 12096
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 9036 12044 9088 12096
rect 10876 12180 10928 12232
rect 11152 12223 11204 12232
rect 11152 12189 11161 12223
rect 11161 12189 11195 12223
rect 11195 12189 11204 12223
rect 11152 12180 11204 12189
rect 11704 12248 11756 12300
rect 15752 12248 15804 12300
rect 16212 12248 16264 12300
rect 16396 12248 16448 12300
rect 19984 12248 20036 12300
rect 23664 12248 23716 12300
rect 25688 12291 25740 12300
rect 25688 12257 25697 12291
rect 25697 12257 25731 12291
rect 25731 12257 25740 12291
rect 25688 12248 25740 12257
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13084 12223 13136 12232
rect 13084 12189 13093 12223
rect 13093 12189 13127 12223
rect 13127 12189 13136 12223
rect 13084 12180 13136 12189
rect 13544 12180 13596 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 16672 12180 16724 12232
rect 17040 12180 17092 12232
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 20352 12180 20404 12232
rect 20720 12180 20772 12232
rect 21640 12180 21692 12232
rect 22008 12223 22060 12232
rect 22008 12189 22017 12223
rect 22017 12189 22051 12223
rect 22051 12189 22060 12223
rect 22008 12180 22060 12189
rect 22284 12223 22336 12232
rect 22284 12189 22293 12223
rect 22293 12189 22327 12223
rect 22327 12189 22336 12223
rect 22284 12180 22336 12189
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 22836 12180 22888 12232
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 25136 12180 25188 12232
rect 26976 12180 27028 12232
rect 28908 12180 28960 12232
rect 11336 12112 11388 12164
rect 14188 12112 14240 12164
rect 13820 12044 13872 12096
rect 14004 12044 14056 12096
rect 14556 12044 14608 12096
rect 17500 12044 17552 12096
rect 17868 12044 17920 12096
rect 19524 12044 19576 12096
rect 23940 12044 23992 12096
rect 24492 12044 24544 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 5632 11840 5684 11892
rect 4068 11772 4120 11824
rect 4804 11772 4856 11824
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 7472 11840 7524 11892
rect 8300 11840 8352 11892
rect 9772 11840 9824 11892
rect 10508 11840 10560 11892
rect 10692 11840 10744 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 7840 11815 7892 11824
rect 7840 11781 7874 11815
rect 7874 11781 7892 11815
rect 7840 11772 7892 11781
rect 8852 11772 8904 11824
rect 10140 11772 10192 11824
rect 7564 11704 7616 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 9128 11704 9180 11756
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 10600 11704 10652 11756
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 7748 11679 7800 11688
rect 7748 11645 7757 11679
rect 7757 11645 7791 11679
rect 7791 11645 7800 11679
rect 7748 11636 7800 11645
rect 5356 11568 5408 11620
rect 7196 11568 7248 11620
rect 9864 11636 9916 11688
rect 8024 11611 8076 11620
rect 8024 11577 8033 11611
rect 8033 11577 8067 11611
rect 8067 11577 8076 11611
rect 8024 11568 8076 11577
rect 8944 11568 8996 11620
rect 9312 11568 9364 11620
rect 9680 11568 9732 11620
rect 10692 11568 10744 11620
rect 3424 11500 3476 11552
rect 6276 11500 6328 11552
rect 8208 11543 8260 11552
rect 8208 11509 8217 11543
rect 8217 11509 8251 11543
rect 8251 11509 8260 11543
rect 10968 11704 11020 11756
rect 11704 11747 11756 11756
rect 11704 11713 11708 11747
rect 11708 11713 11742 11747
rect 11742 11713 11756 11747
rect 11704 11704 11756 11713
rect 11244 11568 11296 11620
rect 11980 11704 12032 11756
rect 14556 11815 14608 11824
rect 14556 11781 14565 11815
rect 14565 11781 14599 11815
rect 14599 11781 14608 11815
rect 14556 11772 14608 11781
rect 16488 11772 16540 11824
rect 24216 11772 24268 11824
rect 12900 11747 12952 11756
rect 12900 11713 12909 11747
rect 12909 11713 12943 11747
rect 12943 11713 12952 11747
rect 12900 11704 12952 11713
rect 12992 11704 13044 11756
rect 12716 11636 12768 11688
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 8208 11500 8260 11509
rect 12532 11543 12584 11552
rect 12532 11509 12541 11543
rect 12541 11509 12575 11543
rect 12575 11509 12584 11543
rect 12532 11500 12584 11509
rect 12900 11500 12952 11552
rect 12992 11500 13044 11552
rect 13544 11704 13596 11756
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 14188 11747 14240 11756
rect 14188 11713 14197 11747
rect 14197 11713 14231 11747
rect 14231 11713 14240 11747
rect 14188 11704 14240 11713
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 17316 11704 17368 11756
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 20720 11704 20772 11756
rect 26424 11704 26476 11756
rect 26884 11704 26936 11756
rect 27988 11840 28040 11892
rect 27528 11747 27580 11756
rect 27528 11713 27537 11747
rect 27537 11713 27571 11747
rect 27571 11713 27580 11747
rect 27528 11704 27580 11713
rect 29000 11704 29052 11756
rect 13728 11568 13780 11620
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 20536 11679 20588 11688
rect 20536 11645 20545 11679
rect 20545 11645 20579 11679
rect 20579 11645 20588 11679
rect 20536 11636 20588 11645
rect 20628 11636 20680 11688
rect 21272 11636 21324 11688
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 27620 11679 27672 11688
rect 27620 11645 27629 11679
rect 27629 11645 27663 11679
rect 27663 11645 27672 11679
rect 27620 11636 27672 11645
rect 15016 11568 15068 11620
rect 21916 11568 21968 11620
rect 14740 11543 14792 11552
rect 14740 11509 14749 11543
rect 14749 11509 14783 11543
rect 14783 11509 14792 11543
rect 14740 11500 14792 11509
rect 19984 11500 20036 11552
rect 21824 11500 21876 11552
rect 23480 11568 23532 11620
rect 22376 11500 22428 11552
rect 23020 11500 23072 11552
rect 24492 11500 24544 11552
rect 28264 11500 28316 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 2228 11296 2280 11348
rect 2596 11296 2648 11348
rect 2688 11296 2740 11348
rect 3424 11296 3476 11348
rect 4988 11296 5040 11348
rect 3148 11228 3200 11280
rect 7564 11296 7616 11348
rect 9128 11296 9180 11348
rect 9312 11296 9364 11348
rect 10600 11339 10652 11348
rect 10600 11305 10609 11339
rect 10609 11305 10643 11339
rect 10643 11305 10652 11339
rect 10600 11296 10652 11305
rect 10692 11296 10744 11348
rect 11520 11296 11572 11348
rect 11612 11339 11664 11348
rect 11612 11305 11621 11339
rect 11621 11305 11655 11339
rect 11655 11305 11664 11339
rect 11612 11296 11664 11305
rect 2688 11135 2740 11144
rect 2688 11101 2697 11135
rect 2697 11101 2731 11135
rect 2731 11101 2740 11135
rect 2688 11092 2740 11101
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 3792 11203 3844 11212
rect 3792 11169 3801 11203
rect 3801 11169 3835 11203
rect 3835 11169 3844 11203
rect 3792 11160 3844 11169
rect 4528 11203 4580 11212
rect 4528 11169 4537 11203
rect 4537 11169 4571 11203
rect 4571 11169 4580 11203
rect 4528 11160 4580 11169
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 3976 11092 4028 11144
rect 9496 11228 9548 11280
rect 10876 11228 10928 11280
rect 11152 11228 11204 11280
rect 6736 11092 6788 11144
rect 8852 11092 8904 11144
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 2964 11024 3016 11076
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 3424 11067 3476 11076
rect 3424 11033 3433 11067
rect 3433 11033 3467 11067
rect 3467 11033 3476 11067
rect 3424 11024 3476 11033
rect 4068 11024 4120 11076
rect 4252 11067 4304 11076
rect 4252 11033 4286 11067
rect 4286 11033 4304 11067
rect 4252 11024 4304 11033
rect 6276 11024 6328 11076
rect 9680 11024 9732 11076
rect 9864 11092 9916 11144
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 10968 11160 11020 11212
rect 12256 11160 12308 11212
rect 11336 11024 11388 11076
rect 11888 11135 11940 11144
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 12900 11160 12952 11212
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 14740 11296 14792 11348
rect 15016 11296 15068 11348
rect 19524 11296 19576 11348
rect 20536 11296 20588 11348
rect 17224 11228 17276 11280
rect 13268 11160 13320 11212
rect 16488 11160 16540 11212
rect 12440 11024 12492 11076
rect 13912 11092 13964 11144
rect 14280 11092 14332 11144
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17868 11092 17920 11144
rect 18512 11092 18564 11144
rect 19064 11092 19116 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 19800 11024 19852 11076
rect 20536 11135 20588 11144
rect 20536 11101 20545 11135
rect 20545 11101 20579 11135
rect 20579 11101 20588 11135
rect 20536 11092 20588 11101
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 20904 11228 20956 11280
rect 22560 11296 22612 11348
rect 23020 11339 23072 11348
rect 23020 11305 23029 11339
rect 23029 11305 23063 11339
rect 23063 11305 23072 11339
rect 23020 11296 23072 11305
rect 27528 11296 27580 11348
rect 29000 11296 29052 11348
rect 21732 11228 21784 11280
rect 21916 11228 21968 11280
rect 22284 11203 22336 11212
rect 22284 11169 22293 11203
rect 22293 11169 22327 11203
rect 22327 11169 22336 11203
rect 22284 11160 22336 11169
rect 22468 11160 22520 11212
rect 22836 11160 22888 11212
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 21272 11067 21324 11076
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 7104 10956 7156 11008
rect 7380 10956 7432 11008
rect 9128 10956 9180 11008
rect 9772 10956 9824 11008
rect 11704 10956 11756 11008
rect 12532 10956 12584 11008
rect 12992 10956 13044 11008
rect 13084 10956 13136 11008
rect 17316 10956 17368 11008
rect 17408 10999 17460 11008
rect 17408 10965 17417 10999
rect 17417 10965 17451 10999
rect 17451 10965 17460 10999
rect 17408 10956 17460 10965
rect 20168 10999 20220 11008
rect 20168 10965 20177 10999
rect 20177 10965 20211 10999
rect 20211 10965 20220 10999
rect 20168 10956 20220 10965
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 21640 11067 21692 11076
rect 21640 11033 21649 11067
rect 21649 11033 21683 11067
rect 21683 11033 21692 11067
rect 21640 11024 21692 11033
rect 23480 11160 23532 11212
rect 24492 11160 24544 11212
rect 27988 11271 28040 11280
rect 27988 11237 27997 11271
rect 27997 11237 28031 11271
rect 28031 11237 28040 11271
rect 27988 11228 28040 11237
rect 21824 11067 21876 11076
rect 21824 11033 21833 11067
rect 21833 11033 21867 11067
rect 21867 11033 21876 11067
rect 21824 11024 21876 11033
rect 26148 11092 26200 11144
rect 26424 11092 26476 11144
rect 27804 11092 27856 11144
rect 28080 11135 28132 11144
rect 28080 11101 28089 11135
rect 28089 11101 28123 11135
rect 28123 11101 28132 11135
rect 28080 11092 28132 11101
rect 28264 11135 28316 11144
rect 28264 11101 28273 11135
rect 28273 11101 28307 11135
rect 28307 11101 28316 11135
rect 28264 11092 28316 11101
rect 28908 11135 28960 11144
rect 28908 11101 28917 11135
rect 28917 11101 28951 11135
rect 28951 11101 28960 11135
rect 28908 11092 28960 11101
rect 29368 11135 29420 11144
rect 29368 11101 29377 11135
rect 29377 11101 29411 11135
rect 29411 11101 29420 11135
rect 29368 11092 29420 11101
rect 23204 11024 23256 11076
rect 25320 10956 25372 11008
rect 27436 11067 27488 11076
rect 27436 11033 27445 11067
rect 27445 11033 27479 11067
rect 27479 11033 27488 11067
rect 27436 11024 27488 11033
rect 26332 10956 26384 11008
rect 27804 10999 27856 11008
rect 27804 10965 27813 10999
rect 27813 10965 27847 10999
rect 27847 10965 27856 10999
rect 27804 10956 27856 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 4252 10752 4304 10804
rect 7196 10752 7248 10804
rect 7748 10752 7800 10804
rect 8944 10752 8996 10804
rect 9772 10752 9824 10804
rect 12900 10752 12952 10804
rect 848 10684 900 10736
rect 2688 10684 2740 10736
rect 6644 10684 6696 10736
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 2872 10616 2924 10668
rect 3976 10659 4028 10668
rect 3976 10625 3985 10659
rect 3985 10625 4019 10659
rect 4019 10625 4028 10659
rect 3976 10616 4028 10625
rect 4528 10616 4580 10668
rect 6552 10616 6604 10668
rect 7104 10616 7156 10668
rect 8852 10684 8904 10736
rect 5724 10591 5776 10600
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9128 10616 9180 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9404 10659 9456 10668
rect 9404 10625 9413 10659
rect 9413 10625 9447 10659
rect 9447 10625 9456 10659
rect 9404 10616 9456 10625
rect 9680 10616 9732 10668
rect 11336 10684 11388 10736
rect 12440 10684 12492 10736
rect 13268 10727 13320 10736
rect 13268 10693 13277 10727
rect 13277 10693 13311 10727
rect 13311 10693 13320 10727
rect 13268 10684 13320 10693
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 9496 10548 9548 10600
rect 10600 10548 10652 10600
rect 10876 10616 10928 10668
rect 13084 10616 13136 10668
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14648 10752 14700 10804
rect 19064 10752 19116 10804
rect 19248 10752 19300 10804
rect 19800 10752 19852 10804
rect 20168 10752 20220 10804
rect 21272 10752 21324 10804
rect 21548 10752 21600 10804
rect 26240 10752 26292 10804
rect 27436 10752 27488 10804
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 14924 10684 14976 10736
rect 17960 10727 18012 10736
rect 15016 10616 15068 10668
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 17960 10693 17969 10727
rect 17969 10693 18003 10727
rect 18003 10693 18012 10727
rect 17960 10684 18012 10693
rect 18420 10684 18472 10736
rect 10968 10548 11020 10600
rect 3240 10480 3292 10532
rect 7196 10480 7248 10532
rect 17040 10548 17092 10600
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17868 10659 17920 10668
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 18880 10616 18932 10668
rect 19708 10616 19760 10668
rect 19984 10684 20036 10736
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 20720 10684 20772 10736
rect 21180 10616 21232 10668
rect 21640 10616 21692 10668
rect 24124 10684 24176 10736
rect 25320 10727 25372 10736
rect 25320 10693 25329 10727
rect 25329 10693 25363 10727
rect 25363 10693 25372 10727
rect 25320 10684 25372 10693
rect 26332 10684 26384 10736
rect 27804 10684 27856 10736
rect 20076 10548 20128 10600
rect 27896 10616 27948 10668
rect 22376 10548 22428 10600
rect 23112 10591 23164 10600
rect 23112 10557 23121 10591
rect 23121 10557 23155 10591
rect 23155 10557 23164 10591
rect 23112 10548 23164 10557
rect 23204 10548 23256 10600
rect 25044 10591 25096 10600
rect 25044 10557 25053 10591
rect 25053 10557 25087 10591
rect 25087 10557 25096 10591
rect 25044 10548 25096 10557
rect 18144 10480 18196 10532
rect 18512 10480 18564 10532
rect 4896 10455 4948 10464
rect 4896 10421 4905 10455
rect 4905 10421 4939 10455
rect 4939 10421 4948 10455
rect 4896 10412 4948 10421
rect 5356 10412 5408 10464
rect 5448 10455 5500 10464
rect 5448 10421 5457 10455
rect 5457 10421 5491 10455
rect 5491 10421 5500 10455
rect 5448 10412 5500 10421
rect 7932 10412 7984 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 8852 10412 8904 10464
rect 9312 10412 9364 10464
rect 10232 10412 10284 10464
rect 10692 10412 10744 10464
rect 11796 10455 11848 10464
rect 11796 10421 11805 10455
rect 11805 10421 11839 10455
rect 11839 10421 11848 10455
rect 11796 10412 11848 10421
rect 12256 10412 12308 10464
rect 13820 10412 13872 10464
rect 17408 10455 17460 10464
rect 17408 10421 17417 10455
rect 17417 10421 17451 10455
rect 17451 10421 17460 10455
rect 17408 10412 17460 10421
rect 18880 10412 18932 10464
rect 19432 10412 19484 10464
rect 21548 10480 21600 10532
rect 28080 10548 28132 10600
rect 20168 10412 20220 10464
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 27988 10455 28040 10464
rect 27988 10421 27997 10455
rect 27997 10421 28031 10455
rect 28031 10421 28040 10455
rect 27988 10412 28040 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3976 10208 4028 10260
rect 5724 10208 5776 10260
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 10508 10208 10560 10260
rect 10876 10208 10928 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 13728 10251 13780 10260
rect 13728 10217 13737 10251
rect 13737 10217 13771 10251
rect 13771 10217 13780 10251
rect 13728 10208 13780 10217
rect 17040 10208 17092 10260
rect 18144 10251 18196 10260
rect 18144 10217 18153 10251
rect 18153 10217 18187 10251
rect 18187 10217 18196 10251
rect 18144 10208 18196 10217
rect 18328 10208 18380 10260
rect 5356 10140 5408 10192
rect 12900 10140 12952 10192
rect 13268 10140 13320 10192
rect 13636 10140 13688 10192
rect 4804 10072 4856 10124
rect 6368 10072 6420 10124
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5448 10004 5500 10056
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8760 10004 8812 10056
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 9956 10047 10008 10056
rect 9956 10013 9965 10047
rect 9965 10013 9999 10047
rect 9999 10013 10008 10047
rect 9956 10004 10008 10013
rect 10048 10004 10100 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 7196 9979 7248 9988
rect 7196 9945 7205 9979
rect 7205 9945 7239 9979
rect 7239 9945 7248 9979
rect 7196 9936 7248 9945
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 10968 10004 11020 10056
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 14280 10072 14332 10124
rect 17500 10072 17552 10124
rect 17868 10140 17920 10192
rect 19340 10208 19392 10260
rect 11796 10004 11848 10013
rect 12624 10004 12676 10056
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 11336 9936 11388 9988
rect 11612 9936 11664 9988
rect 13084 9979 13136 9988
rect 13084 9945 13093 9979
rect 13093 9945 13127 9979
rect 13127 9945 13136 9979
rect 13084 9936 13136 9945
rect 14004 9936 14056 9988
rect 14372 9936 14424 9988
rect 14924 9936 14976 9988
rect 17316 9979 17368 9988
rect 17316 9945 17325 9979
rect 17325 9945 17359 9979
rect 17359 9945 17368 9979
rect 17316 9936 17368 9945
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 4804 9868 4856 9920
rect 7288 9868 7340 9920
rect 10140 9868 10192 9920
rect 17868 9868 17920 9920
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19432 10072 19484 10124
rect 19616 10208 19668 10260
rect 19892 10208 19944 10260
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 23112 10208 23164 10260
rect 24124 10251 24176 10260
rect 24124 10217 24133 10251
rect 24133 10217 24167 10251
rect 24167 10217 24176 10251
rect 24124 10208 24176 10217
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 23204 10072 23256 10124
rect 23664 10072 23716 10124
rect 18420 9979 18472 9988
rect 18420 9945 18429 9979
rect 18429 9945 18463 9979
rect 18463 9945 18472 9979
rect 18420 9936 18472 9945
rect 19708 10004 19760 10056
rect 21732 10047 21784 10056
rect 21732 10013 21741 10047
rect 21741 10013 21775 10047
rect 21775 10013 21784 10047
rect 21732 10004 21784 10013
rect 26424 10208 26476 10260
rect 27896 10208 27948 10260
rect 26332 10115 26384 10124
rect 26332 10081 26341 10115
rect 26341 10081 26375 10115
rect 26375 10081 26384 10115
rect 26332 10072 26384 10081
rect 26240 10004 26292 10056
rect 27620 10115 27672 10124
rect 27620 10081 27629 10115
rect 27629 10081 27663 10115
rect 27663 10081 27672 10115
rect 27620 10072 27672 10081
rect 27988 10072 28040 10124
rect 29000 10004 29052 10056
rect 27620 9936 27672 9988
rect 27804 9868 27856 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4804 9664 4856 9716
rect 9036 9664 9088 9716
rect 10048 9664 10100 9716
rect 10968 9664 11020 9716
rect 11428 9664 11480 9716
rect 2136 9596 2188 9648
rect 4528 9596 4580 9648
rect 6000 9596 6052 9648
rect 7196 9596 7248 9648
rect 4160 9528 4212 9580
rect 6736 9528 6788 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 9404 9639 9456 9648
rect 9404 9605 9421 9639
rect 9421 9605 9456 9639
rect 9404 9596 9456 9605
rect 9220 9571 9272 9580
rect 11612 9596 11664 9648
rect 13728 9707 13780 9716
rect 13728 9673 13737 9707
rect 13737 9673 13771 9707
rect 13771 9673 13780 9707
rect 13728 9664 13780 9673
rect 17500 9664 17552 9716
rect 18420 9664 18472 9716
rect 20904 9664 20956 9716
rect 13268 9596 13320 9648
rect 14924 9639 14976 9648
rect 14924 9605 14933 9639
rect 14933 9605 14967 9639
rect 14967 9605 14976 9639
rect 14924 9596 14976 9605
rect 21640 9664 21692 9716
rect 1308 9460 1360 9512
rect 2320 9460 2372 9512
rect 2688 9460 2740 9512
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4712 9460 4764 9512
rect 6828 9392 6880 9444
rect 2688 9324 2740 9376
rect 4620 9324 4672 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7012 9324 7064 9376
rect 9220 9537 9262 9571
rect 9262 9537 9272 9571
rect 9220 9528 9272 9537
rect 8852 9460 8904 9512
rect 9496 9460 9548 9512
rect 9588 9460 9640 9512
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 13544 9528 13596 9580
rect 11888 9460 11940 9512
rect 13084 9460 13136 9512
rect 13728 9528 13780 9580
rect 16672 9528 16724 9580
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 20260 9528 20312 9580
rect 19248 9460 19300 9512
rect 9588 9324 9640 9376
rect 10232 9392 10284 9444
rect 12992 9392 13044 9444
rect 21180 9528 21232 9580
rect 22100 9596 22152 9648
rect 22928 9596 22980 9648
rect 23756 9596 23808 9648
rect 24216 9596 24268 9648
rect 26332 9596 26384 9648
rect 27344 9596 27396 9648
rect 29000 9639 29052 9648
rect 29000 9605 29009 9639
rect 29009 9605 29043 9639
rect 29043 9605 29052 9639
rect 29000 9596 29052 9605
rect 21548 9528 21600 9580
rect 21916 9460 21968 9512
rect 23572 9571 23624 9580
rect 23572 9537 23581 9571
rect 23581 9537 23615 9571
rect 23615 9537 23624 9571
rect 23572 9528 23624 9537
rect 24124 9528 24176 9580
rect 28908 9528 28960 9580
rect 23664 9460 23716 9512
rect 25044 9460 25096 9512
rect 27712 9460 27764 9512
rect 21088 9392 21140 9444
rect 11888 9324 11940 9376
rect 12164 9367 12216 9376
rect 12164 9333 12173 9367
rect 12173 9333 12207 9367
rect 12207 9333 12216 9367
rect 12164 9324 12216 9333
rect 15568 9324 15620 9376
rect 17592 9324 17644 9376
rect 18972 9324 19024 9376
rect 26884 9392 26936 9444
rect 23388 9324 23440 9376
rect 24860 9324 24912 9376
rect 29368 9435 29420 9444
rect 29368 9401 29377 9435
rect 29377 9401 29411 9435
rect 29411 9401 29420 9435
rect 29368 9392 29420 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 2320 9163 2372 9172
rect 2320 9129 2329 9163
rect 2329 9129 2363 9163
rect 2363 9129 2372 9163
rect 2320 9120 2372 9129
rect 6736 9120 6788 9172
rect 7564 9120 7616 9172
rect 9680 9120 9732 9172
rect 10232 9120 10284 9172
rect 2596 8984 2648 9036
rect 3148 8984 3200 9036
rect 4620 8984 4672 9036
rect 2320 8916 2372 8968
rect 2504 8916 2556 8968
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 2688 8916 2740 8925
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 5264 8848 5316 8900
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 8852 8984 8904 9036
rect 9036 8984 9088 9036
rect 9588 8984 9640 9036
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 6000 8848 6052 8857
rect 6460 8780 6512 8832
rect 7104 8848 7156 8900
rect 7196 8891 7248 8900
rect 7196 8857 7205 8891
rect 7205 8857 7239 8891
rect 7239 8857 7248 8891
rect 7196 8848 7248 8857
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 10508 8959 10560 8968
rect 10508 8925 10517 8959
rect 10517 8925 10551 8959
rect 10551 8925 10560 8959
rect 10508 8916 10560 8925
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 11796 8916 11848 8968
rect 11244 8848 11296 8900
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 12900 8959 12952 8968
rect 12900 8925 12909 8959
rect 12909 8925 12943 8959
rect 12943 8925 12952 8959
rect 12900 8916 12952 8925
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 13176 9120 13228 9172
rect 16948 9163 17000 9172
rect 16948 9129 16957 9163
rect 16957 9129 16991 9163
rect 16991 9129 17000 9163
rect 16948 9120 17000 9129
rect 15660 8984 15712 9036
rect 16396 8984 16448 9036
rect 10232 8823 10284 8832
rect 10232 8789 10241 8823
rect 10241 8789 10275 8823
rect 10275 8789 10284 8823
rect 10232 8780 10284 8789
rect 10508 8780 10560 8832
rect 15568 8959 15620 8968
rect 15568 8925 15577 8959
rect 15577 8925 15611 8959
rect 15611 8925 15620 8959
rect 15568 8916 15620 8925
rect 17040 8916 17092 8968
rect 22008 9120 22060 9172
rect 22100 9120 22152 9172
rect 27344 9163 27396 9172
rect 27344 9129 27353 9163
rect 27353 9129 27387 9163
rect 27387 9129 27396 9163
rect 27344 9120 27396 9129
rect 19248 9095 19300 9104
rect 19248 9061 19257 9095
rect 19257 9061 19291 9095
rect 19291 9061 19300 9095
rect 19248 9052 19300 9061
rect 22192 9052 22244 9104
rect 20720 8984 20772 9036
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 17592 8959 17644 8968
rect 17592 8925 17601 8959
rect 17601 8925 17635 8959
rect 17635 8925 17644 8959
rect 17592 8916 17644 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 21088 8959 21140 8968
rect 21088 8925 21097 8959
rect 21097 8925 21131 8959
rect 21131 8925 21140 8959
rect 23112 8984 23164 9036
rect 21088 8916 21140 8925
rect 22376 8916 22428 8968
rect 23388 8959 23440 8968
rect 23388 8925 23397 8959
rect 23397 8925 23431 8959
rect 23431 8925 23440 8959
rect 23388 8916 23440 8925
rect 23480 8959 23532 8968
rect 23480 8925 23525 8959
rect 23525 8925 23532 8959
rect 23480 8916 23532 8925
rect 11888 8780 11940 8832
rect 20076 8848 20128 8900
rect 23296 8891 23348 8900
rect 14740 8780 14792 8832
rect 16212 8780 16264 8832
rect 16672 8780 16724 8832
rect 17684 8780 17736 8832
rect 18236 8823 18288 8832
rect 18236 8789 18245 8823
rect 18245 8789 18279 8823
rect 18279 8789 18288 8823
rect 18236 8780 18288 8789
rect 19708 8780 19760 8832
rect 23296 8857 23305 8891
rect 23305 8857 23339 8891
rect 23339 8857 23348 8891
rect 23296 8848 23348 8857
rect 24492 8959 24544 8968
rect 24492 8925 24501 8959
rect 24501 8925 24535 8959
rect 24535 8925 24544 8959
rect 24492 8916 24544 8925
rect 26424 8916 26476 8968
rect 20904 8780 20956 8832
rect 23848 8848 23900 8900
rect 28632 8848 28684 8900
rect 23572 8780 23624 8832
rect 24676 8780 24728 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5264 8576 5316 8628
rect 7196 8576 7248 8628
rect 9128 8576 9180 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 12808 8576 12860 8628
rect 13820 8576 13872 8628
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 7564 8551 7616 8560
rect 7564 8517 7573 8551
rect 7573 8517 7607 8551
rect 7607 8517 7616 8551
rect 7564 8508 7616 8517
rect 11244 8508 11296 8560
rect 14740 8551 14792 8560
rect 14740 8517 14749 8551
rect 14749 8517 14783 8551
rect 14783 8517 14792 8551
rect 14740 8508 14792 8517
rect 15476 8508 15528 8560
rect 16120 8508 16172 8560
rect 2320 8440 2372 8492
rect 5632 8440 5684 8492
rect 6920 8440 6972 8492
rect 12348 8440 12400 8492
rect 12440 8440 12492 8492
rect 12992 8440 13044 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 6828 8372 6880 8424
rect 7472 8415 7524 8424
rect 7472 8381 7481 8415
rect 7481 8381 7515 8415
rect 7515 8381 7524 8415
rect 7472 8372 7524 8381
rect 9404 8372 9456 8424
rect 12532 8372 12584 8424
rect 13452 8372 13504 8424
rect 13728 8372 13780 8424
rect 14280 8440 14332 8492
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17868 8576 17920 8628
rect 18236 8576 18288 8628
rect 19708 8576 19760 8628
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 23480 8576 23532 8628
rect 23664 8576 23716 8628
rect 24124 8619 24176 8628
rect 24124 8585 24133 8619
rect 24133 8585 24167 8619
rect 24167 8585 24176 8619
rect 24124 8576 24176 8585
rect 24952 8576 25004 8628
rect 26884 8576 26936 8628
rect 17040 8440 17092 8492
rect 17224 8440 17276 8492
rect 17684 8508 17736 8560
rect 17592 8440 17644 8492
rect 19248 8440 19300 8492
rect 22192 8508 22244 8560
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20352 8483 20404 8492
rect 20352 8449 20362 8483
rect 20362 8449 20396 8483
rect 20396 8449 20404 8483
rect 20352 8440 20404 8449
rect 20628 8440 20680 8492
rect 2412 8304 2464 8356
rect 16396 8372 16448 8424
rect 23480 8440 23532 8492
rect 23664 8483 23716 8492
rect 23664 8449 23673 8483
rect 23673 8449 23707 8483
rect 23707 8449 23716 8483
rect 23664 8440 23716 8449
rect 23296 8372 23348 8424
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 28172 8440 28224 8492
rect 29276 8483 29328 8492
rect 29276 8449 29285 8483
rect 29285 8449 29319 8483
rect 29319 8449 29328 8483
rect 29276 8440 29328 8449
rect 23848 8347 23900 8356
rect 23848 8313 23857 8347
rect 23857 8313 23891 8347
rect 23891 8313 23900 8347
rect 23848 8304 23900 8313
rect 24124 8304 24176 8356
rect 1768 8236 1820 8288
rect 8024 8236 8076 8288
rect 9864 8236 9916 8288
rect 10968 8236 11020 8288
rect 11612 8236 11664 8288
rect 12440 8236 12492 8288
rect 20536 8236 20588 8288
rect 20904 8236 20956 8288
rect 21916 8236 21968 8288
rect 23388 8236 23440 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 7288 8032 7340 8084
rect 10324 8075 10376 8084
rect 10324 8041 10333 8075
rect 10333 8041 10367 8075
rect 10367 8041 10376 8075
rect 10324 8032 10376 8041
rect 11704 8032 11756 8084
rect 12624 8032 12676 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 15476 8032 15528 8084
rect 21272 8032 21324 8084
rect 22284 8032 22336 8084
rect 4712 7964 4764 7973
rect 848 7828 900 7880
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 4804 7896 4856 7948
rect 5816 7896 5868 7948
rect 5908 7939 5960 7948
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 9404 7964 9456 8016
rect 10968 8007 11020 8016
rect 10968 7973 10977 8007
rect 10977 7973 11011 8007
rect 11011 7973 11020 8007
rect 10968 7964 11020 7973
rect 11060 7964 11112 8016
rect 5724 7828 5776 7880
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 4436 7760 4488 7812
rect 6368 7760 6420 7812
rect 7288 7828 7340 7880
rect 8024 7828 8076 7880
rect 6000 7692 6052 7744
rect 7564 7760 7616 7812
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 9496 7828 9548 7880
rect 10048 7828 10100 7880
rect 10324 7828 10376 7880
rect 8484 7760 8536 7812
rect 10416 7760 10468 7812
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11704 7896 11756 7948
rect 11796 7828 11848 7880
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 13820 7896 13872 7948
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 13912 7828 13964 7880
rect 14188 7828 14240 7880
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 16672 7828 16724 7880
rect 18052 7828 18104 7880
rect 19248 7828 19300 7880
rect 19340 7828 19392 7880
rect 19892 7896 19944 7948
rect 20168 7896 20220 7948
rect 20076 7828 20128 7880
rect 20628 7896 20680 7948
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7104 7692 7156 7744
rect 7932 7692 7984 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 12072 7803 12124 7812
rect 12072 7769 12081 7803
rect 12081 7769 12115 7803
rect 12115 7769 12124 7803
rect 12072 7760 12124 7769
rect 12164 7760 12216 7812
rect 19984 7760 20036 7812
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 20996 7939 21048 7948
rect 20996 7905 21005 7939
rect 21005 7905 21039 7939
rect 21039 7905 21048 7939
rect 20996 7896 21048 7905
rect 21824 8007 21876 8016
rect 21824 7973 21833 8007
rect 21833 7973 21867 8007
rect 21867 7973 21876 8007
rect 21824 7964 21876 7973
rect 22652 7964 22704 8016
rect 22836 8032 22888 8084
rect 24032 8032 24084 8084
rect 24124 8032 24176 8084
rect 11060 7692 11112 7744
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 17684 7692 17736 7744
rect 19432 7692 19484 7744
rect 20168 7735 20220 7744
rect 20168 7701 20177 7735
rect 20177 7701 20211 7735
rect 20211 7701 20220 7735
rect 20168 7692 20220 7701
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 22560 7896 22612 7948
rect 22100 7828 22152 7880
rect 22284 7871 22336 7880
rect 22284 7837 22288 7871
rect 22288 7837 22322 7871
rect 22322 7837 22336 7871
rect 22284 7828 22336 7837
rect 22376 7871 22428 7880
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 22652 7871 22704 7880
rect 22652 7837 22660 7871
rect 22660 7837 22694 7871
rect 22694 7837 22704 7871
rect 22652 7828 22704 7837
rect 22744 7871 22796 7880
rect 22744 7837 22753 7871
rect 22753 7837 22787 7871
rect 22787 7837 22796 7871
rect 22744 7828 22796 7837
rect 21456 7803 21508 7812
rect 21456 7769 21465 7803
rect 21465 7769 21499 7803
rect 21499 7769 21508 7803
rect 21456 7760 21508 7769
rect 21548 7803 21600 7812
rect 21548 7769 21557 7803
rect 21557 7769 21591 7803
rect 21591 7769 21600 7803
rect 21548 7760 21600 7769
rect 22100 7735 22152 7744
rect 22100 7701 22109 7735
rect 22109 7701 22143 7735
rect 22143 7701 22152 7735
rect 22100 7692 22152 7701
rect 22284 7692 22336 7744
rect 22560 7760 22612 7812
rect 23204 7828 23256 7880
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 23480 7828 23532 7837
rect 23848 7760 23900 7812
rect 24216 7871 24268 7880
rect 24216 7837 24225 7871
rect 24225 7837 24259 7871
rect 24259 7837 24268 7871
rect 24216 7828 24268 7837
rect 24400 7828 24452 7880
rect 29552 7896 29604 7948
rect 24676 7871 24728 7880
rect 24676 7837 24685 7871
rect 24685 7837 24719 7871
rect 24719 7837 24728 7871
rect 24676 7828 24728 7837
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 29368 7871 29420 7880
rect 29368 7837 29377 7871
rect 29377 7837 29411 7871
rect 29411 7837 29420 7871
rect 29368 7828 29420 7837
rect 24308 7760 24360 7812
rect 29736 7760 29788 7812
rect 29184 7735 29236 7744
rect 29184 7701 29193 7735
rect 29193 7701 29227 7735
rect 29227 7701 29236 7735
rect 29184 7692 29236 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 6552 7488 6604 7540
rect 8208 7488 8260 7540
rect 8300 7488 8352 7540
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 1676 7148 1728 7200
rect 4436 7259 4488 7268
rect 4436 7225 4445 7259
rect 4445 7225 4479 7259
rect 4479 7225 4488 7259
rect 4436 7216 4488 7225
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 6092 7420 6144 7472
rect 7288 7420 7340 7472
rect 5724 7352 5776 7361
rect 6184 7352 6236 7404
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 6644 7284 6696 7336
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 6000 7216 6052 7268
rect 6552 7216 6604 7268
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 8576 7395 8628 7404
rect 8576 7361 8585 7395
rect 8585 7361 8619 7395
rect 8619 7361 8628 7395
rect 8576 7352 8628 7361
rect 10416 7488 10468 7540
rect 11520 7488 11572 7540
rect 12716 7488 12768 7540
rect 12900 7488 12952 7540
rect 13084 7488 13136 7540
rect 14372 7488 14424 7540
rect 15660 7488 15712 7540
rect 17960 7488 18012 7540
rect 19708 7488 19760 7540
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 20628 7488 20680 7540
rect 9128 7284 9180 7336
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 10232 7352 10284 7404
rect 10876 7420 10928 7472
rect 11060 7352 11112 7404
rect 12624 7420 12676 7472
rect 11244 7352 11296 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 9864 7284 9916 7336
rect 10508 7259 10560 7268
rect 10508 7225 10517 7259
rect 10517 7225 10551 7259
rect 10551 7225 10560 7259
rect 10508 7216 10560 7225
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 11428 7216 11480 7268
rect 11980 7352 12032 7404
rect 12348 7352 12400 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 13544 7352 13596 7404
rect 12440 7284 12492 7336
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 13728 7284 13780 7336
rect 14004 7352 14056 7404
rect 14648 7420 14700 7472
rect 14464 7352 14516 7404
rect 16580 7352 16632 7404
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 17684 7395 17736 7404
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 17960 7395 18012 7404
rect 17960 7361 17969 7395
rect 17969 7361 18003 7395
rect 18003 7361 18012 7395
rect 17960 7352 18012 7361
rect 19892 7420 19944 7472
rect 18052 7284 18104 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 19708 7395 19760 7404
rect 19708 7361 19717 7395
rect 19717 7361 19751 7395
rect 19751 7361 19760 7395
rect 19708 7352 19760 7361
rect 19524 7284 19576 7336
rect 20076 7352 20128 7404
rect 20904 7420 20956 7472
rect 22100 7488 22152 7540
rect 22284 7488 22336 7540
rect 22652 7488 22704 7540
rect 24216 7488 24268 7540
rect 21548 7420 21600 7472
rect 21916 7420 21968 7472
rect 20996 7352 21048 7404
rect 21456 7395 21508 7404
rect 21456 7361 21465 7395
rect 21465 7361 21499 7395
rect 21499 7361 21508 7395
rect 21456 7352 21508 7361
rect 21824 7352 21876 7404
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 23296 7352 23348 7404
rect 24676 7420 24728 7472
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 23112 7284 23164 7336
rect 23848 7284 23900 7336
rect 24584 7284 24636 7336
rect 29828 7284 29880 7336
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10968 7148 11020 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 17500 7148 17552 7200
rect 19708 7148 19760 7200
rect 21180 7148 21232 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1676 6987 1728 6996
rect 1676 6953 1706 6987
rect 1706 6953 1728 6987
rect 1676 6944 1728 6953
rect 2964 6944 3016 6996
rect 7748 6944 7800 6996
rect 8576 6944 8628 6996
rect 10232 6944 10284 6996
rect 12808 6944 12860 6996
rect 15292 6987 15344 6996
rect 15292 6953 15301 6987
rect 15301 6953 15335 6987
rect 15335 6953 15344 6987
rect 15292 6944 15344 6953
rect 17960 6944 18012 6996
rect 18604 6944 18656 6996
rect 18696 6944 18748 6996
rect 6828 6876 6880 6928
rect 9772 6876 9824 6928
rect 1308 6808 1360 6860
rect 4068 6808 4120 6860
rect 4620 6808 4672 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 4712 6740 4764 6792
rect 8392 6808 8444 6860
rect 12348 6808 12400 6860
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 8484 6740 8536 6792
rect 2412 6672 2464 6724
rect 4804 6647 4856 6656
rect 4804 6613 4813 6647
rect 4813 6613 4847 6647
rect 4847 6613 4856 6647
rect 4804 6604 4856 6613
rect 9220 6740 9272 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10968 6740 11020 6792
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 11796 6672 11848 6724
rect 12348 6715 12400 6724
rect 12348 6681 12357 6715
rect 12357 6681 12391 6715
rect 12391 6681 12400 6715
rect 12348 6672 12400 6681
rect 12716 6808 12768 6860
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 12624 6740 12676 6792
rect 13268 6740 13320 6792
rect 15016 6808 15068 6860
rect 11704 6604 11756 6656
rect 15292 6672 15344 6724
rect 15568 6783 15620 6792
rect 15568 6749 15577 6783
rect 15577 6749 15611 6783
rect 15611 6749 15620 6783
rect 15568 6740 15620 6749
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 16764 6808 16816 6860
rect 17224 6808 17276 6860
rect 16120 6740 16172 6792
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 17960 6808 18012 6860
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 19524 6808 19576 6860
rect 19708 6808 19760 6860
rect 19248 6740 19300 6792
rect 20076 6876 20128 6928
rect 16672 6672 16724 6724
rect 14096 6604 14148 6656
rect 15200 6604 15252 6656
rect 15660 6604 15712 6656
rect 17592 6672 17644 6724
rect 19892 6740 19944 6792
rect 17224 6604 17276 6656
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 19340 6604 19392 6656
rect 19616 6715 19668 6724
rect 19616 6681 19625 6715
rect 19625 6681 19659 6715
rect 19659 6681 19668 6715
rect 19616 6672 19668 6681
rect 19708 6672 19760 6724
rect 23940 6672 23992 6724
rect 20168 6604 20220 6656
rect 21088 6647 21140 6656
rect 21088 6613 21097 6647
rect 21097 6613 21131 6647
rect 21131 6613 21140 6647
rect 21088 6604 21140 6613
rect 21364 6604 21416 6656
rect 29092 6604 29144 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 8208 6400 8260 6452
rect 848 6264 900 6316
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 8484 6400 8536 6452
rect 9128 6400 9180 6452
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 12900 6400 12952 6452
rect 10416 6332 10468 6384
rect 11796 6375 11848 6384
rect 11796 6341 11805 6375
rect 11805 6341 11839 6375
rect 11839 6341 11848 6375
rect 11796 6332 11848 6341
rect 11888 6375 11940 6384
rect 11888 6341 11897 6375
rect 11897 6341 11931 6375
rect 11931 6341 11940 6375
rect 11888 6332 11940 6341
rect 6644 6239 6696 6248
rect 6644 6205 6653 6239
rect 6653 6205 6687 6239
rect 6687 6205 6696 6239
rect 6644 6196 6696 6205
rect 8576 6264 8628 6316
rect 9496 6264 9548 6316
rect 9128 6196 9180 6248
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 11152 6264 11204 6316
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 10968 6196 11020 6248
rect 11060 6196 11112 6248
rect 12072 6307 12124 6316
rect 12072 6273 12081 6307
rect 12081 6273 12115 6307
rect 12115 6273 12124 6307
rect 12072 6264 12124 6273
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 13912 6307 13964 6316
rect 13912 6273 13921 6307
rect 13921 6273 13955 6307
rect 13955 6273 13964 6307
rect 13912 6264 13964 6273
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 7012 6128 7064 6180
rect 8760 6128 8812 6180
rect 15384 6196 15436 6248
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 17316 6400 17368 6452
rect 20260 6400 20312 6452
rect 17132 6375 17184 6384
rect 17132 6341 17141 6375
rect 17141 6341 17175 6375
rect 17175 6341 17184 6375
rect 17132 6332 17184 6341
rect 17224 6375 17276 6384
rect 17224 6341 17233 6375
rect 17233 6341 17267 6375
rect 17267 6341 17276 6375
rect 17224 6332 17276 6341
rect 17592 6332 17644 6384
rect 18236 6332 18288 6384
rect 19432 6264 19484 6316
rect 19892 6264 19944 6316
rect 19708 6196 19760 6248
rect 19800 6196 19852 6248
rect 20444 6264 20496 6316
rect 21640 6332 21692 6384
rect 21456 6307 21508 6316
rect 21456 6273 21464 6307
rect 21464 6273 21498 6307
rect 21498 6273 21508 6307
rect 21456 6264 21508 6273
rect 21548 6307 21600 6316
rect 21548 6273 21557 6307
rect 21557 6273 21591 6307
rect 21591 6273 21600 6307
rect 21548 6264 21600 6273
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 21180 6196 21232 6248
rect 22560 6264 22612 6316
rect 24492 6400 24544 6452
rect 22836 6307 22888 6316
rect 22836 6273 22845 6307
rect 22845 6273 22879 6307
rect 22879 6273 22888 6307
rect 22836 6264 22888 6273
rect 17132 6128 17184 6180
rect 20260 6128 20312 6180
rect 10232 6060 10284 6112
rect 11704 6060 11756 6112
rect 11796 6060 11848 6112
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 17040 6060 17092 6112
rect 18236 6060 18288 6112
rect 20168 6060 20220 6112
rect 23204 6264 23256 6316
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 23756 6264 23808 6316
rect 23848 6307 23900 6316
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 24124 6307 24176 6316
rect 24124 6273 24133 6307
rect 24133 6273 24167 6307
rect 24167 6273 24176 6307
rect 24124 6264 24176 6273
rect 24308 6307 24360 6316
rect 24308 6273 24317 6307
rect 24317 6273 24351 6307
rect 24351 6273 24360 6307
rect 24308 6264 24360 6273
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 29092 6307 29144 6316
rect 29092 6273 29101 6307
rect 29101 6273 29135 6307
rect 29135 6273 29144 6307
rect 29092 6264 29144 6273
rect 23940 6128 23992 6180
rect 29368 6239 29420 6248
rect 29368 6205 29377 6239
rect 29377 6205 29411 6239
rect 29411 6205 29420 6239
rect 29368 6196 29420 6205
rect 24584 6128 24636 6180
rect 24768 6060 24820 6112
rect 24952 6060 25004 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 10140 5856 10192 5908
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 11520 5899 11572 5908
rect 11520 5865 11529 5899
rect 11529 5865 11563 5899
rect 11563 5865 11572 5899
rect 11520 5856 11572 5865
rect 13820 5856 13872 5908
rect 13912 5856 13964 5908
rect 16488 5856 16540 5908
rect 8576 5788 8628 5840
rect 11060 5788 11112 5840
rect 3148 5720 3200 5772
rect 5448 5720 5500 5772
rect 7472 5720 7524 5772
rect 8760 5763 8812 5772
rect 8760 5729 8769 5763
rect 8769 5729 8803 5763
rect 8803 5729 8812 5763
rect 8760 5720 8812 5729
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 5540 5652 5592 5704
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7380 5652 7432 5704
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8944 5652 8996 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 11612 5720 11664 5772
rect 15476 5788 15528 5840
rect 16672 5856 16724 5908
rect 17316 5856 17368 5908
rect 17408 5856 17460 5908
rect 18512 5856 18564 5908
rect 19248 5856 19300 5908
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 9220 5652 9272 5661
rect 4436 5627 4488 5636
rect 4436 5593 4445 5627
rect 4445 5593 4479 5627
rect 4479 5593 4488 5627
rect 4436 5584 4488 5593
rect 8852 5584 8904 5636
rect 10324 5695 10376 5704
rect 9588 5584 9640 5636
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 12624 5652 12676 5704
rect 13084 5695 13136 5704
rect 13084 5661 13091 5695
rect 13091 5661 13136 5695
rect 13084 5652 13136 5661
rect 13452 5652 13504 5704
rect 13820 5652 13872 5704
rect 14648 5695 14700 5704
rect 14648 5661 14657 5695
rect 14657 5661 14691 5695
rect 14691 5661 14700 5695
rect 14648 5652 14700 5661
rect 15752 5652 15804 5704
rect 5908 5559 5960 5568
rect 5908 5525 5917 5559
rect 5917 5525 5951 5559
rect 5951 5525 5960 5559
rect 5908 5516 5960 5525
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 10140 5516 10192 5568
rect 13176 5627 13228 5636
rect 13176 5593 13185 5627
rect 13185 5593 13219 5627
rect 13219 5593 13228 5627
rect 13176 5584 13228 5593
rect 13268 5627 13320 5636
rect 13268 5593 13277 5627
rect 13277 5593 13311 5627
rect 13311 5593 13320 5627
rect 13268 5584 13320 5593
rect 15660 5584 15712 5636
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 18604 5788 18656 5840
rect 21548 5788 21600 5840
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 29644 5788 29696 5840
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17224 5695 17276 5704
rect 17224 5661 17233 5695
rect 17233 5661 17267 5695
rect 17267 5661 17276 5695
rect 17224 5652 17276 5661
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 17684 5652 17736 5704
rect 17500 5627 17552 5636
rect 17500 5593 17509 5627
rect 17509 5593 17543 5627
rect 17543 5593 17552 5627
rect 17500 5584 17552 5593
rect 21824 5720 21876 5772
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 19064 5652 19116 5704
rect 19524 5652 19576 5704
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 20444 5652 20496 5704
rect 19248 5584 19300 5636
rect 21088 5695 21140 5704
rect 21088 5661 21097 5695
rect 21097 5661 21131 5695
rect 21131 5661 21140 5695
rect 21088 5652 21140 5661
rect 21364 5695 21416 5704
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 23756 5720 23808 5772
rect 21364 5652 21416 5661
rect 22928 5695 22980 5704
rect 22928 5661 22937 5695
rect 22937 5661 22971 5695
rect 22971 5661 22980 5695
rect 22928 5652 22980 5661
rect 23848 5652 23900 5704
rect 21456 5584 21508 5636
rect 24584 5695 24636 5704
rect 24584 5661 24593 5695
rect 24593 5661 24627 5695
rect 24627 5661 24636 5695
rect 24584 5652 24636 5661
rect 24768 5695 24820 5704
rect 24768 5661 24777 5695
rect 24777 5661 24811 5695
rect 24811 5661 24820 5695
rect 24768 5652 24820 5661
rect 24952 5695 25004 5704
rect 24952 5661 24961 5695
rect 24961 5661 24995 5695
rect 24995 5661 25004 5695
rect 24952 5652 25004 5661
rect 19708 5516 19760 5568
rect 20076 5516 20128 5568
rect 20996 5516 21048 5568
rect 21272 5516 21324 5568
rect 21640 5516 21692 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4436 5312 4488 5364
rect 4804 5312 4856 5364
rect 5540 5312 5592 5364
rect 8024 5312 8076 5364
rect 8484 5312 8536 5364
rect 9956 5312 10008 5364
rect 11980 5312 12032 5364
rect 13820 5312 13872 5364
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 14648 5312 14700 5364
rect 16488 5355 16540 5364
rect 16488 5321 16497 5355
rect 16497 5321 16531 5355
rect 16531 5321 16540 5355
rect 16488 5312 16540 5321
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 20168 5312 20220 5364
rect 22192 5312 22244 5364
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 5908 5244 5960 5296
rect 6644 5287 6696 5296
rect 6644 5253 6653 5287
rect 6653 5253 6687 5287
rect 6687 5253 6696 5287
rect 6644 5244 6696 5253
rect 8576 5244 8628 5296
rect 848 5176 900 5228
rect 4160 5176 4212 5228
rect 5448 5108 5500 5160
rect 5632 5176 5684 5228
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9220 5176 9272 5228
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10692 5176 10744 5228
rect 11060 5219 11112 5228
rect 11060 5185 11069 5219
rect 11069 5185 11103 5219
rect 11103 5185 11112 5219
rect 11060 5176 11112 5185
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 11612 5176 11664 5228
rect 11980 5176 12032 5228
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 18604 5287 18656 5296
rect 18604 5253 18613 5287
rect 18613 5253 18647 5287
rect 18647 5253 18656 5287
rect 18604 5244 18656 5253
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 13820 5176 13872 5228
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 14832 5176 14884 5228
rect 15108 5219 15160 5228
rect 15108 5185 15117 5219
rect 15117 5185 15151 5219
rect 15151 5185 15160 5219
rect 15108 5176 15160 5185
rect 5632 5040 5684 5092
rect 13452 5108 13504 5160
rect 14004 5108 14056 5160
rect 15016 5108 15068 5160
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15568 5176 15620 5228
rect 16120 5219 16172 5228
rect 16120 5185 16129 5219
rect 16129 5185 16163 5219
rect 16163 5185 16172 5219
rect 16120 5176 16172 5185
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 16764 5176 16816 5228
rect 17224 5176 17276 5228
rect 17316 5219 17368 5228
rect 17316 5185 17325 5219
rect 17325 5185 17359 5219
rect 17359 5185 17368 5219
rect 17316 5176 17368 5185
rect 17408 5219 17460 5228
rect 17408 5185 17417 5219
rect 17417 5185 17451 5219
rect 17451 5185 17460 5219
rect 17408 5176 17460 5185
rect 17592 5176 17644 5228
rect 9036 5040 9088 5092
rect 9128 5040 9180 5092
rect 11244 5040 11296 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 11888 4972 11940 5024
rect 13084 5040 13136 5092
rect 15384 5083 15436 5092
rect 15384 5049 15393 5083
rect 15393 5049 15427 5083
rect 15427 5049 15436 5083
rect 15384 5040 15436 5049
rect 16120 5040 16172 5092
rect 17224 5040 17276 5092
rect 18512 5176 18564 5228
rect 18972 5176 19024 5228
rect 19340 5176 19392 5228
rect 19524 5219 19576 5228
rect 19524 5185 19533 5219
rect 19533 5185 19567 5219
rect 19567 5185 19576 5219
rect 19524 5176 19576 5185
rect 20076 5219 20128 5228
rect 20076 5185 20085 5219
rect 20085 5185 20119 5219
rect 20119 5185 20128 5219
rect 20076 5176 20128 5185
rect 21272 5176 21324 5228
rect 22284 5176 22336 5228
rect 22468 5219 22520 5228
rect 22468 5185 22477 5219
rect 22477 5185 22511 5219
rect 22511 5185 22520 5219
rect 22468 5176 22520 5185
rect 22652 5219 22704 5228
rect 22652 5185 22660 5219
rect 22660 5185 22694 5219
rect 22694 5185 22704 5219
rect 22652 5176 22704 5185
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 23848 5176 23900 5228
rect 29276 5219 29328 5228
rect 29276 5185 29285 5219
rect 29285 5185 29319 5219
rect 29319 5185 29328 5219
rect 29276 5176 29328 5185
rect 17040 4972 17092 5024
rect 17132 4972 17184 5024
rect 18972 5040 19024 5092
rect 19064 5083 19116 5092
rect 19064 5049 19073 5083
rect 19073 5049 19107 5083
rect 19107 5049 19116 5083
rect 19064 5040 19116 5049
rect 18788 4972 18840 5024
rect 21088 4972 21140 5024
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 8852 4768 8904 4820
rect 13084 4768 13136 4820
rect 1584 4700 1636 4752
rect 10048 4700 10100 4752
rect 10140 4700 10192 4752
rect 12072 4700 12124 4752
rect 14372 4768 14424 4820
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 14924 4768 14976 4820
rect 15568 4768 15620 4820
rect 16580 4768 16632 4820
rect 17408 4768 17460 4820
rect 18512 4811 18564 4820
rect 18512 4777 18521 4811
rect 18521 4777 18555 4811
rect 18555 4777 18564 4811
rect 18512 4768 18564 4777
rect 22744 4768 22796 4820
rect 17132 4700 17184 4752
rect 17316 4700 17368 4752
rect 19432 4700 19484 4752
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 11888 4607 11940 4616
rect 11888 4573 11897 4607
rect 11897 4573 11931 4607
rect 11931 4573 11940 4607
rect 11888 4564 11940 4573
rect 12624 4564 12676 4616
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 13268 4607 13320 4616
rect 13268 4573 13277 4607
rect 13277 4573 13311 4607
rect 13311 4573 13320 4607
rect 13268 4564 13320 4573
rect 13544 4632 13596 4684
rect 14740 4564 14792 4616
rect 11980 4496 12032 4548
rect 12256 4496 12308 4548
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 15476 4564 15528 4616
rect 16672 4564 16724 4616
rect 16856 4564 16908 4616
rect 19248 4632 19300 4684
rect 21916 4675 21968 4684
rect 21916 4641 21925 4675
rect 21925 4641 21959 4675
rect 21959 4641 21968 4675
rect 22468 4743 22520 4752
rect 22468 4709 22477 4743
rect 22477 4709 22511 4743
rect 22511 4709 22520 4743
rect 22468 4700 22520 4709
rect 22652 4700 22704 4752
rect 21916 4632 21968 4641
rect 17684 4496 17736 4548
rect 11060 4428 11112 4480
rect 11612 4428 11664 4480
rect 17316 4428 17368 4480
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 19432 4564 19484 4616
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 24124 4768 24176 4820
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 23112 4607 23164 4616
rect 23112 4573 23151 4607
rect 23151 4573 23164 4607
rect 23112 4564 23164 4573
rect 23480 4564 23532 4616
rect 21180 4496 21232 4548
rect 20444 4471 20496 4480
rect 20444 4437 20453 4471
rect 20453 4437 20487 4471
rect 20487 4437 20496 4471
rect 20444 4428 20496 4437
rect 23204 4428 23256 4480
rect 23664 4564 23716 4616
rect 24124 4564 24176 4616
rect 25320 4564 25372 4616
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 24492 4428 24544 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 9956 4156 10008 4208
rect 10968 4199 11020 4208
rect 10968 4165 10977 4199
rect 10977 4165 11011 4199
rect 11011 4165 11020 4199
rect 11888 4224 11940 4276
rect 10968 4156 11020 4165
rect 6368 4088 6420 4140
rect 11244 4156 11296 4208
rect 11796 4088 11848 4140
rect 12256 4156 12308 4208
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 13268 4224 13320 4276
rect 15476 4224 15528 4276
rect 17224 4224 17276 4276
rect 19064 4224 19116 4276
rect 19248 4224 19300 4276
rect 20352 4224 20404 4276
rect 25320 4224 25372 4276
rect 12624 4156 12676 4208
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 13820 4156 13872 4208
rect 14556 4156 14608 4208
rect 13452 4088 13504 4140
rect 14832 4088 14884 4140
rect 13636 4020 13688 4072
rect 13176 3952 13228 4004
rect 14648 3952 14700 4004
rect 16396 4020 16448 4072
rect 17592 4088 17644 4140
rect 20444 4156 20496 4208
rect 23756 4199 23808 4208
rect 23756 4165 23765 4199
rect 23765 4165 23799 4199
rect 23799 4165 23808 4199
rect 23756 4156 23808 4165
rect 24492 4156 24544 4208
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 18236 4088 18288 4140
rect 17960 3952 18012 4004
rect 13360 3884 13412 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 16580 3884 16632 3936
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 19708 4063 19760 4072
rect 19708 4029 19717 4063
rect 19717 4029 19751 4063
rect 19751 4029 19760 4063
rect 19708 4020 19760 4029
rect 23296 4020 23348 4072
rect 20720 3884 20772 3936
rect 21088 3884 21140 3936
rect 22560 3884 22612 3936
rect 22652 3884 22704 3936
rect 22928 3884 22980 3936
rect 23388 3884 23440 3936
rect 24124 4020 24176 4072
rect 25044 3884 25096 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 11060 3680 11112 3732
rect 12716 3723 12768 3732
rect 12716 3689 12725 3723
rect 12725 3689 12759 3723
rect 12759 3689 12768 3723
rect 12716 3680 12768 3689
rect 13268 3680 13320 3732
rect 13636 3723 13688 3732
rect 13636 3689 13645 3723
rect 13645 3689 13679 3723
rect 13679 3689 13688 3723
rect 13636 3680 13688 3689
rect 16580 3723 16632 3732
rect 16580 3689 16589 3723
rect 16589 3689 16623 3723
rect 16623 3689 16632 3723
rect 16580 3680 16632 3689
rect 17960 3723 18012 3732
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 18052 3680 18104 3732
rect 10968 3612 11020 3664
rect 16672 3612 16724 3664
rect 17868 3612 17920 3664
rect 18420 3655 18472 3664
rect 18420 3621 18429 3655
rect 18429 3621 18463 3655
rect 18463 3621 18472 3655
rect 18420 3612 18472 3621
rect 11244 3544 11296 3596
rect 848 3476 900 3528
rect 9036 3476 9088 3528
rect 9588 3476 9640 3528
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11152 3408 11204 3460
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 11980 3408 12032 3460
rect 14280 3544 14332 3596
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15292 3544 15344 3596
rect 19340 3544 19392 3596
rect 13084 3476 13136 3528
rect 13452 3476 13504 3528
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 19708 3612 19760 3664
rect 22284 3612 22336 3664
rect 22468 3655 22520 3664
rect 22468 3621 22477 3655
rect 22477 3621 22511 3655
rect 22511 3621 22520 3655
rect 22468 3612 22520 3621
rect 22560 3655 22612 3664
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 23112 3723 23164 3732
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 23388 3680 23440 3732
rect 23664 3680 23716 3732
rect 21088 3544 21140 3596
rect 22744 3544 22796 3596
rect 23388 3544 23440 3596
rect 13820 3451 13872 3460
rect 13820 3417 13829 3451
rect 13829 3417 13863 3451
rect 13863 3417 13872 3451
rect 13820 3408 13872 3417
rect 15384 3408 15436 3460
rect 16856 3408 16908 3460
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 16396 3340 16448 3392
rect 17592 3383 17644 3392
rect 17592 3349 17601 3383
rect 17601 3349 17635 3383
rect 17635 3349 17644 3383
rect 17592 3340 17644 3349
rect 18144 3408 18196 3460
rect 20720 3519 20772 3528
rect 20720 3485 20729 3519
rect 20729 3485 20763 3519
rect 20763 3485 20772 3519
rect 20720 3476 20772 3485
rect 22468 3476 22520 3528
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 23756 3519 23808 3528
rect 23756 3485 23765 3519
rect 23765 3485 23799 3519
rect 23799 3485 23808 3519
rect 23756 3476 23808 3485
rect 20352 3408 20404 3460
rect 20628 3451 20680 3460
rect 20628 3417 20637 3451
rect 20637 3417 20671 3451
rect 20671 3417 20680 3451
rect 20628 3408 20680 3417
rect 18604 3340 18656 3392
rect 19708 3340 19760 3392
rect 21272 3408 21324 3460
rect 22008 3408 22060 3460
rect 22468 3340 22520 3392
rect 22836 3383 22888 3392
rect 22836 3349 22845 3383
rect 22845 3349 22879 3383
rect 22879 3349 22888 3383
rect 22836 3340 22888 3349
rect 23480 3340 23532 3392
rect 24124 3476 24176 3528
rect 29276 3451 29328 3460
rect 29276 3417 29285 3451
rect 29285 3417 29319 3451
rect 29319 3417 29328 3451
rect 29276 3408 29328 3417
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1860 3136 1912 3188
rect 11336 3136 11388 3188
rect 11980 3136 12032 3188
rect 12164 3136 12216 3188
rect 664 2932 716 2984
rect 11704 3068 11756 3120
rect 14280 3136 14332 3188
rect 14740 3136 14792 3188
rect 9588 3000 9640 3052
rect 11612 2932 11664 2984
rect 848 2864 900 2916
rect 1584 2796 1636 2848
rect 11520 2864 11572 2916
rect 12072 3000 12124 3052
rect 13268 3111 13320 3120
rect 13268 3077 13277 3111
rect 13277 3077 13311 3111
rect 13311 3077 13320 3111
rect 13268 3068 13320 3077
rect 15384 3136 15436 3188
rect 16120 3111 16172 3120
rect 16120 3077 16129 3111
rect 16129 3077 16163 3111
rect 16163 3077 16172 3111
rect 16120 3068 16172 3077
rect 16672 3068 16724 3120
rect 17868 3068 17920 3120
rect 16488 3000 16540 3052
rect 17040 3000 17092 3052
rect 19340 3068 19392 3120
rect 19708 3068 19760 3120
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 22008 3136 22060 3188
rect 22928 3136 22980 3188
rect 20720 3068 20772 3120
rect 17592 2932 17644 2984
rect 18144 2932 18196 2984
rect 19432 2932 19484 2984
rect 22560 3043 22612 3052
rect 22560 3009 22569 3043
rect 22569 3009 22603 3043
rect 22603 3009 22612 3043
rect 22560 3000 22612 3009
rect 22744 3043 22796 3052
rect 22744 3009 22753 3043
rect 22753 3009 22787 3043
rect 22787 3009 22796 3043
rect 22744 3000 22796 3009
rect 23756 3136 23808 3188
rect 20628 2932 20680 2984
rect 23480 3068 23532 3120
rect 28724 3111 28776 3120
rect 28724 3077 28733 3111
rect 28733 3077 28767 3111
rect 28767 3077 28776 3111
rect 28724 3068 28776 3077
rect 23296 3043 23348 3052
rect 23296 3009 23305 3043
rect 23305 3009 23339 3043
rect 23339 3009 23348 3043
rect 23296 3000 23348 3009
rect 25320 3043 25372 3052
rect 25320 3009 25329 3043
rect 25329 3009 25363 3043
rect 25363 3009 25372 3043
rect 25320 3000 25372 3009
rect 29000 3000 29052 3052
rect 29368 3000 29420 3052
rect 23572 2975 23624 2984
rect 23572 2941 23581 2975
rect 23581 2941 23615 2975
rect 23615 2941 23624 2975
rect 23572 2932 23624 2941
rect 11888 2796 11940 2848
rect 11980 2796 12032 2848
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 22008 2864 22060 2916
rect 20352 2796 20404 2848
rect 22928 2864 22980 2916
rect 29092 2907 29144 2916
rect 29092 2873 29101 2907
rect 29101 2873 29135 2907
rect 29135 2873 29144 2907
rect 29092 2864 29144 2873
rect 23388 2796 23440 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 8208 2592 8260 2644
rect 8668 2592 8720 2644
rect 10416 2592 10468 2644
rect 12072 2592 12124 2644
rect 12808 2592 12860 2644
rect 16212 2635 16264 2644
rect 16212 2601 16221 2635
rect 16221 2601 16255 2635
rect 16255 2601 16264 2635
rect 16212 2592 16264 2601
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 4988 2567 5040 2576
rect 4988 2533 4997 2567
rect 4997 2533 5031 2567
rect 5031 2533 5040 2567
rect 4988 2524 5040 2533
rect 19524 2592 19576 2644
rect 23112 2592 23164 2644
rect 23296 2592 23348 2644
rect 23572 2635 23624 2644
rect 23572 2601 23581 2635
rect 23581 2601 23615 2635
rect 23615 2601 23624 2635
rect 23572 2592 23624 2601
rect 23664 2635 23716 2644
rect 23664 2601 23673 2635
rect 23673 2601 23707 2635
rect 23707 2601 23716 2635
rect 23664 2592 23716 2601
rect 17684 2524 17736 2576
rect 21180 2524 21232 2576
rect 940 2388 992 2440
rect 1952 2388 2004 2440
rect 3240 2388 3292 2440
rect 20 2320 72 2372
rect 4528 2320 4580 2372
rect 5816 2388 5868 2440
rect 7104 2388 7156 2440
rect 7748 2388 7800 2440
rect 8300 2456 8352 2508
rect 10140 2456 10192 2508
rect 10600 2456 10652 2508
rect 8852 2388 8904 2440
rect 9036 2388 9088 2440
rect 10324 2388 10376 2440
rect 11888 2456 11940 2508
rect 23664 2456 23716 2508
rect 8944 2320 8996 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 8024 2252 8076 2304
rect 12808 2388 12860 2440
rect 12900 2388 12952 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 11612 2320 11664 2372
rect 14188 2320 14240 2372
rect 15476 2320 15528 2372
rect 16120 2388 16172 2440
rect 16488 2388 16540 2440
rect 16580 2320 16632 2372
rect 17408 2388 17460 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19984 2388 20036 2440
rect 22560 2388 22612 2440
rect 23296 2388 23348 2440
rect 24492 2388 24544 2440
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 18696 2320 18748 2372
rect 19340 2363 19392 2372
rect 19340 2329 19349 2363
rect 19349 2329 19383 2363
rect 19383 2329 19392 2363
rect 19340 2320 19392 2329
rect 23112 2320 23164 2372
rect 23388 2363 23440 2372
rect 23388 2329 23413 2363
rect 23413 2329 23440 2363
rect 23388 2320 23440 2329
rect 25780 2320 25832 2372
rect 15568 2252 15620 2304
rect 15660 2252 15712 2304
rect 18880 2295 18932 2304
rect 18880 2261 18889 2295
rect 18889 2261 18923 2295
rect 18923 2261 18932 2295
rect 18880 2252 18932 2261
rect 20812 2252 20864 2304
rect 27068 2320 27120 2372
rect 27252 2295 27304 2304
rect 27252 2261 27261 2295
rect 27261 2261 27295 2295
rect 27295 2261 27304 2295
rect 27252 2252 27304 2261
rect 28172 2295 28224 2304
rect 28172 2261 28181 2295
rect 28181 2261 28215 2295
rect 28215 2261 28224 2295
rect 28172 2252 28224 2261
rect 28356 2320 28408 2372
rect 29644 2388 29696 2440
rect 29276 2363 29328 2372
rect 29276 2329 29285 2363
rect 29285 2329 29319 2363
rect 29319 2329 29328 2363
rect 29276 2320 29328 2329
rect 29184 2295 29236 2304
rect 29184 2261 29193 2295
rect 29193 2261 29227 2295
rect 29227 2261 29236 2295
rect 29184 2252 29236 2261
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 14004 1980 14056 2032
rect 28172 1980 28224 2032
rect 1584 1912 1636 1964
rect 21916 1912 21968 1964
rect 13268 1844 13320 1896
rect 19616 1844 19668 1896
rect 11428 1776 11480 1828
rect 27252 1776 27304 1828
rect 14464 1640 14516 1692
rect 29184 1640 29236 1692
<< metal2 >>
rect 18 32247 74 33047
rect 938 32736 994 32745
rect 938 32671 994 32680
rect 32 30258 60 32247
rect 20 30252 72 30258
rect 20 30194 72 30200
rect 848 30184 900 30190
rect 846 30152 848 30161
rect 900 30152 902 30161
rect 846 30087 902 30096
rect 952 29714 980 32671
rect 1306 32247 1362 33047
rect 2594 32247 2650 33047
rect 3882 32247 3938 33047
rect 5170 32247 5226 33047
rect 6458 32247 6514 33047
rect 7102 32247 7158 33047
rect 8390 32247 8446 33047
rect 9678 32247 9734 33047
rect 10966 32247 11022 33047
rect 12254 32247 12310 33047
rect 13542 32247 13598 33047
rect 14830 32247 14886 33047
rect 15474 32247 15530 33047
rect 16762 32247 16818 33047
rect 18050 32247 18106 33047
rect 19338 32247 19394 33047
rect 20626 32247 20682 33047
rect 21914 32247 21970 33047
rect 22558 32247 22614 33047
rect 23846 32247 23902 33047
rect 25134 32247 25190 33047
rect 26422 32247 26478 33047
rect 27710 32247 27766 33047
rect 28998 32247 29054 33047
rect 29366 32736 29422 32745
rect 29366 32671 29422 32680
rect 1214 31376 1270 31385
rect 1214 31311 1270 31320
rect 940 29708 992 29714
rect 940 29650 992 29656
rect 1228 29578 1256 31311
rect 1320 30326 1348 32247
rect 2608 30326 2636 32247
rect 1308 30320 1360 30326
rect 1308 30262 1360 30268
rect 2596 30320 2648 30326
rect 2596 30262 2648 30268
rect 3896 30258 3924 32247
rect 5184 31226 5212 32247
rect 5184 31198 5304 31226
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5276 30258 5304 31198
rect 7116 30258 7144 32247
rect 8404 30326 8432 32247
rect 9692 30326 9720 32247
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 9680 30320 9732 30326
rect 9680 30262 9732 30268
rect 10980 30258 11008 32247
rect 12268 30258 12296 32247
rect 13556 30258 13584 32247
rect 14844 30258 14872 32247
rect 15488 30326 15516 32247
rect 15476 30320 15528 30326
rect 15476 30262 15528 30268
rect 16776 30258 16804 32247
rect 18064 30258 18092 32247
rect 19352 30326 19380 32247
rect 20640 30326 20668 32247
rect 21928 30326 21956 32247
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 22572 30258 22600 32247
rect 23860 30258 23888 32247
rect 25148 30326 25176 32247
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 26436 30258 26464 32247
rect 27724 30326 27752 32247
rect 28538 31376 28594 31385
rect 28538 31311 28594 31320
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 3884 30252 3936 30258
rect 3884 30194 3936 30200
rect 5264 30252 5316 30258
rect 5264 30194 5316 30200
rect 7104 30252 7156 30258
rect 7104 30194 7156 30200
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 13544 30252 13596 30258
rect 13544 30194 13596 30200
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 16764 30252 16816 30258
rect 16764 30194 16816 30200
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 23848 30252 23900 30258
rect 23848 30194 23900 30200
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 1952 30184 2004 30190
rect 1952 30126 2004 30132
rect 11612 30184 11664 30190
rect 11612 30126 11664 30132
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 1216 29572 1268 29578
rect 1216 29514 1268 29520
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28665 1440 29106
rect 1398 28656 1454 28665
rect 1398 28591 1454 28600
rect 848 27464 900 27470
rect 846 27432 848 27441
rect 1676 27464 1728 27470
rect 900 27432 902 27441
rect 1676 27406 1728 27412
rect 846 27367 902 27376
rect 1492 26308 1544 26314
rect 1492 26250 1544 26256
rect 1504 25945 1532 26250
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 848 24812 900 24818
rect 848 24754 900 24760
rect 860 24721 888 24754
rect 846 24712 902 24721
rect 846 24647 902 24656
rect 846 23760 902 23769
rect 846 23695 848 23704
rect 900 23695 902 23704
rect 848 23666 900 23672
rect 848 22568 900 22574
rect 848 22510 900 22516
rect 860 22409 888 22510
rect 846 22400 902 22409
rect 846 22335 902 22344
rect 1688 22001 1716 27406
rect 1674 21992 1730 22001
rect 1674 21927 1730 21936
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 860 21321 888 21490
rect 1768 21412 1820 21418
rect 1768 21354 1820 21360
rect 846 21312 902 21321
rect 846 21247 902 21256
rect 1400 20868 1452 20874
rect 1400 20810 1452 20816
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 1412 19378 1440 20810
rect 1676 19848 1728 19854
rect 1674 19816 1676 19825
rect 1728 19816 1730 19825
rect 1674 19751 1730 19760
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19446 1716 19654
rect 1676 19440 1728 19446
rect 1676 19382 1728 19388
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 848 18760 900 18766
rect 848 18702 900 18708
rect 860 18601 888 18702
rect 846 18592 902 18601
rect 846 18527 902 18536
rect 848 17264 900 17270
rect 846 17232 848 17241
rect 900 17232 902 17241
rect 846 17167 902 17176
rect 848 16584 900 16590
rect 846 16552 848 16561
rect 900 16552 902 16561
rect 846 16487 902 16496
rect 1584 16516 1636 16522
rect 1584 16458 1636 16464
rect 1596 15706 1624 16458
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 1504 15065 1532 15370
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 848 12232 900 12238
rect 846 12200 848 12209
rect 900 12200 902 12209
rect 846 12135 902 12144
rect 846 10840 902 10849
rect 846 10775 902 10784
rect 860 10742 888 10775
rect 848 10736 900 10742
rect 848 10678 900 10684
rect 1674 10704 1730 10713
rect 1674 10639 1676 10648
rect 1728 10639 1730 10648
rect 1676 10610 1728 10616
rect 1308 9512 1360 9518
rect 1308 9454 1360 9460
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1320 6866 1348 9454
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1780 8294 1808 21354
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1768 8288 1820 8294
rect 1398 8256 1454 8265
rect 1768 8230 1820 8236
rect 1398 8191 1454 8200
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 7002 1716 7142
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1308 6860 1360 6866
rect 1308 6802 1360 6808
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 1584 5024 1636 5030
rect 846 4992 902 5001
rect 1584 4966 1636 4972
rect 846 4927 902 4936
rect 1596 4758 1624 4966
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 846 3632 902 3641
rect 846 3567 902 3576
rect 860 3534 888 3567
rect 848 3528 900 3534
rect 848 3470 900 3476
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 676 800 704 2926
rect 848 2916 900 2922
rect 848 2858 900 2864
rect 860 921 888 2858
rect 1596 2854 1624 3334
rect 1872 3194 1900 18226
rect 1964 14890 1992 30126
rect 2688 30116 2740 30122
rect 2688 30058 2740 30064
rect 2964 30116 3016 30122
rect 2964 30058 3016 30064
rect 3332 30116 3384 30122
rect 3332 30058 3384 30064
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 2596 29572 2648 29578
rect 2596 29514 2648 29520
rect 2044 26308 2096 26314
rect 2044 26250 2096 26256
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 12918 1992 13806
rect 1952 12912 2004 12918
rect 1952 12854 2004 12860
rect 1952 12164 2004 12170
rect 1952 12106 2004 12112
rect 1964 5817 1992 12106
rect 2056 7993 2084 26250
rect 2608 26042 2636 29514
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 2148 17882 2176 18226
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12918 2176 13126
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2228 12096 2280 12102
rect 2228 12038 2280 12044
rect 2240 11354 2268 12038
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2148 9178 2176 9590
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2332 9178 2360 9454
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2332 8498 2360 8910
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2042 7984 2098 7993
rect 2042 7919 2098 7928
rect 2332 6322 2360 8434
rect 2424 8362 2452 24550
rect 2700 23050 2728 30058
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2688 23044 2740 23050
rect 2688 22986 2740 22992
rect 2686 22672 2742 22681
rect 2792 22642 2820 24210
rect 2686 22607 2688 22616
rect 2740 22607 2742 22616
rect 2780 22636 2832 22642
rect 2688 22578 2740 22584
rect 2780 22578 2832 22584
rect 2792 21554 2820 22578
rect 2976 22166 3004 30058
rect 3344 26858 3372 30058
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 5448 30048 5500 30054
rect 5448 29990 5500 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4712 29096 4764 29102
rect 4712 29038 4764 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4724 28082 4752 29038
rect 5276 28762 5304 29990
rect 5264 28756 5316 28762
rect 5264 28698 5316 28704
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4712 28076 4764 28082
rect 4712 28018 4764 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3700 27532 3752 27538
rect 3700 27474 3752 27480
rect 3332 26852 3384 26858
rect 3332 26794 3384 26800
rect 3712 25906 3740 27474
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4724 26382 4752 28018
rect 4802 27568 4858 27577
rect 4802 27503 4804 27512
rect 4856 27503 4858 27512
rect 4804 27474 4856 27480
rect 5356 27396 5408 27402
rect 5356 27338 5408 27344
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5368 27130 5396 27338
rect 5356 27124 5408 27130
rect 5356 27066 5408 27072
rect 5460 26602 5488 29990
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7564 28552 7616 28558
rect 7564 28494 7616 28500
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 7300 28218 7328 28494
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 6552 28076 6604 28082
rect 6552 28018 6604 28024
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5828 27402 5856 27814
rect 5816 27396 5868 27402
rect 5816 27338 5868 27344
rect 5368 26574 5488 26602
rect 4804 26444 4856 26450
rect 4804 26386 4856 26392
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4160 26308 4212 26314
rect 4160 26250 4212 26256
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3712 24274 3740 25842
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3988 25498 4016 25774
rect 4172 25684 4200 26250
rect 4620 26240 4672 26246
rect 4620 26182 4672 26188
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4080 25656 4200 25684
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 4080 25242 4108 25656
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25498 4660 26182
rect 4724 25974 4752 26182
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 3988 25214 4108 25242
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 3884 25152 3936 25158
rect 3884 25094 3936 25100
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3252 23866 3280 24142
rect 3896 24070 3924 25094
rect 3884 24064 3936 24070
rect 3884 24006 3936 24012
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 3068 22234 3096 22510
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 3896 21894 3924 24006
rect 3988 23730 4016 25214
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4252 24336 4304 24342
rect 4252 24278 4304 24284
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4172 23730 4200 24210
rect 4264 23866 4292 24278
rect 4620 24268 4672 24274
rect 4620 24210 4672 24216
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4344 24064 4396 24070
rect 4344 24006 4396 24012
rect 4252 23860 4304 23866
rect 4252 23802 4304 23808
rect 4356 23730 4384 24006
rect 4540 23798 4568 24142
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4344 23724 4396 23730
rect 4344 23666 4396 23672
rect 3988 21944 4016 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 24210
rect 4724 23526 4752 25230
rect 4816 24342 4844 26386
rect 5368 26330 5396 26574
rect 5264 26308 5316 26314
rect 5368 26302 5488 26330
rect 5264 26250 5316 26256
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5172 24948 5224 24954
rect 5172 24890 5224 24896
rect 5184 24342 5212 24890
rect 5276 24682 5304 26250
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5368 26042 5396 26182
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5368 24954 5396 25978
rect 5356 24948 5408 24954
rect 5356 24890 5408 24896
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 5368 24410 5396 24754
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 5172 24336 5224 24342
rect 5172 24278 5224 24284
rect 5184 24052 5212 24278
rect 5184 24024 5304 24052
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4804 23860 4856 23866
rect 4804 23802 4856 23808
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4448 22778 4476 23122
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4160 22636 4212 22642
rect 4160 22578 4212 22584
rect 4172 22420 4200 22578
rect 4080 22392 4200 22420
rect 4080 22098 4108 22392
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 22234 4660 23258
rect 4816 23118 4844 23802
rect 5276 23798 5304 24024
rect 5264 23792 5316 23798
rect 5264 23734 5316 23740
rect 4896 23724 4948 23730
rect 4896 23666 4948 23672
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 4816 22710 4844 23054
rect 4908 22982 4936 23666
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5368 23118 5396 23598
rect 5356 23112 5408 23118
rect 5354 23080 5356 23089
rect 5408 23080 5410 23089
rect 5264 23044 5316 23050
rect 5354 23015 5410 23024
rect 5264 22986 5316 22992
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4068 21956 4120 21962
rect 3988 21916 4068 21944
rect 4068 21898 4120 21904
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3884 21616 3936 21622
rect 3884 21558 3936 21564
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2792 20874 2820 21490
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2596 19712 2648 19718
rect 2596 19654 2648 19660
rect 2608 18426 2636 19654
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2792 18970 2820 19314
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2884 18766 2912 19790
rect 3160 18970 3188 21422
rect 3896 21146 3924 21558
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 4080 20942 4108 21898
rect 4724 21894 4752 22374
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3528 20466 3556 20810
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3424 19780 3476 19786
rect 3424 19722 3476 19728
rect 3436 19446 3464 19722
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2516 17678 2544 17818
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2884 16658 2912 18702
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3160 17610 3188 18226
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3344 17678 3372 18158
rect 3436 17882 3464 19382
rect 3804 19378 3832 20334
rect 4080 19854 4108 20878
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3884 18692 3936 18698
rect 3884 18634 3936 18640
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 3344 17338 3372 17614
rect 3436 17610 3464 17818
rect 3792 17672 3844 17678
rect 3792 17614 3844 17620
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2596 16176 2648 16182
rect 2596 16118 2648 16124
rect 2608 15706 2636 16118
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2884 15502 2912 16594
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15502 3372 16050
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3620 15706 3648 15982
rect 3712 15706 3740 17206
rect 3804 17202 3832 17614
rect 3896 17542 3924 18634
rect 4080 17882 4108 18702
rect 4172 18290 4200 18770
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4264 18154 4292 18770
rect 4356 18698 4384 18906
rect 4632 18698 4660 21422
rect 4816 20618 4844 22646
rect 5276 22234 5304 22986
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5356 21956 5408 21962
rect 5356 21898 5408 21904
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4724 20590 4844 20618
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4448 18426 4476 18634
rect 4436 18420 4488 18426
rect 4436 18362 4488 18368
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4172 17678 4200 17750
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4264 17542 4292 17614
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3804 15502 3832 16118
rect 3896 16114 3924 17478
rect 4356 17202 4384 17682
rect 4528 17332 4580 17338
rect 4632 17320 4660 18226
rect 4580 17292 4660 17320
rect 4528 17274 4580 17280
rect 4724 17218 4752 20590
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4816 20058 4844 20470
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4896 19984 4948 19990
rect 4816 19932 4896 19938
rect 4816 19926 4948 19932
rect 4816 19910 4936 19926
rect 4816 19394 4844 19910
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4816 19366 4936 19394
rect 4908 19310 4936 19366
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4908 18970 4936 19246
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 5092 18902 5120 19314
rect 5080 18896 5132 18902
rect 5080 18838 5132 18844
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4816 17746 4844 18702
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4344 17196 4396 17202
rect 4724 17190 4844 17218
rect 4344 17138 4396 17144
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16114 4660 17002
rect 4724 16182 4752 17070
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 4252 16108 4304 16114
rect 4620 16108 4672 16114
rect 4304 16068 4620 16096
rect 4252 16050 4304 16056
rect 4620 16050 4672 16056
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15502 4016 15914
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4080 15502 4108 15642
rect 4632 15502 4660 15846
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 2516 14396 2544 15438
rect 2780 14408 2832 14414
rect 2516 14368 2780 14396
rect 2516 13326 2544 14368
rect 2780 14350 2832 14356
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12442 2544 13262
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2516 8974 2544 12378
rect 2608 11354 2636 13330
rect 3344 12374 3372 15438
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 14006 3464 14214
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13530 3832 13670
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3528 12986 3556 13262
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3436 12238 3464 12718
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2700 11234 2728 11290
rect 3160 11286 3188 12174
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3436 11354 3464 11494
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 2608 11206 2728 11234
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2608 10674 2636 11206
rect 3160 11150 3188 11222
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 2700 10742 2728 11086
rect 3436 11082 3464 11290
rect 3804 11218 3832 12922
rect 3988 12782 4016 15438
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4080 13870 4108 15098
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4816 14634 4844 17190
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15570 5212 16050
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4632 14606 4844 14634
rect 4632 13938 4660 14606
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13326 4108 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4080 12850 4108 13262
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12776 4028 12782
rect 4028 12724 4108 12730
rect 3976 12718 4108 12724
rect 3988 12702 4108 12718
rect 4080 12306 4108 12702
rect 4632 12646 4660 13874
rect 4724 13870 4752 14282
rect 4816 14074 4844 14418
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12374 4752 13330
rect 4816 12918 4844 14010
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3988 11150 4016 12242
rect 4080 11830 4108 12242
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4080 11082 4108 11766
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2872 10668 2924 10674
rect 2976 10656 3004 11018
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 2924 10628 3004 10656
rect 2872 10610 2924 10616
rect 2608 9602 2636 10610
rect 3252 10538 3280 10950
rect 4264 10810 4292 11018
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3988 10266 4016 10610
rect 4264 10554 4292 10746
rect 4540 10674 4568 11154
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4080 10526 4292 10554
rect 3976 10260 4028 10266
rect 4080 10248 4108 10526
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10220 4200 10248
rect 3976 10202 4028 10208
rect 2608 9574 2728 9602
rect 2608 9042 2636 9574
rect 2700 9518 2728 9574
rect 3988 9518 4016 10202
rect 4172 9586 4200 10220
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9654 4568 9862
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4724 9518 4752 12310
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4816 11218 4844 11766
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11354 5028 11698
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4816 10130 4844 11154
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 10062 4936 10406
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9722 4844 9862
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 5276 9674 5304 18226
rect 5368 18154 5396 21898
rect 5460 18290 5488 26302
rect 5724 25900 5776 25906
rect 5724 25842 5776 25848
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5644 24682 5672 24890
rect 5736 24818 5764 25842
rect 5920 25294 5948 28018
rect 6460 27872 6512 27878
rect 6460 27814 6512 27820
rect 6368 27600 6420 27606
rect 6368 27542 6420 27548
rect 6380 27402 6408 27542
rect 6472 27470 6500 27814
rect 6564 27606 6592 28018
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 6552 27600 6604 27606
rect 6552 27542 6604 27548
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6828 27464 6880 27470
rect 7116 27441 7144 27950
rect 6828 27406 6880 27412
rect 7102 27432 7158 27441
rect 6368 27396 6420 27402
rect 6368 27338 6420 27344
rect 6184 27056 6236 27062
rect 6184 26998 6236 27004
rect 6000 26308 6052 26314
rect 6000 26250 6052 26256
rect 6012 26042 6040 26250
rect 6000 26036 6052 26042
rect 6000 25978 6052 25984
rect 6012 25294 6040 25978
rect 6092 25968 6144 25974
rect 6092 25910 6144 25916
rect 5908 25288 5960 25294
rect 5908 25230 5960 25236
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 5908 24948 5960 24954
rect 5908 24890 5960 24896
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 5632 24676 5684 24682
rect 5632 24618 5684 24624
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5552 24206 5580 24346
rect 5540 24200 5592 24206
rect 5540 24142 5592 24148
rect 5644 23322 5672 24618
rect 5920 24206 5948 24890
rect 6104 24614 6132 25910
rect 6196 25158 6224 26998
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6288 25906 6316 26182
rect 6276 25900 6328 25906
rect 6276 25842 6328 25848
rect 6276 25424 6328 25430
rect 6276 25366 6328 25372
rect 6184 25152 6236 25158
rect 6184 25094 6236 25100
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 6012 23526 6040 24006
rect 6104 23730 6132 24550
rect 6288 24410 6316 25366
rect 6380 25294 6408 27338
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6656 27130 6684 27270
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6840 27062 6868 27406
rect 7102 27367 7104 27376
rect 7156 27367 7158 27376
rect 7104 27338 7156 27344
rect 7300 27062 7328 28154
rect 7484 27946 7512 28358
rect 7472 27940 7524 27946
rect 7472 27882 7524 27888
rect 7484 27470 7512 27882
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 6840 26790 6868 26998
rect 6920 26988 6972 26994
rect 6920 26930 6972 26936
rect 6932 26790 6960 26930
rect 7392 26926 7420 27406
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7392 26790 7420 26862
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6920 26784 6972 26790
rect 6920 26726 6972 26732
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 6644 26376 6696 26382
rect 6644 26318 6696 26324
rect 6460 26240 6512 26246
rect 6460 26182 6512 26188
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6184 24268 6236 24274
rect 6288 24256 6316 24346
rect 6236 24228 6316 24256
rect 6184 24210 6236 24216
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 6000 23520 6052 23526
rect 6000 23462 6052 23468
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5540 23044 5592 23050
rect 5540 22986 5592 22992
rect 5552 22710 5580 22986
rect 5540 22704 5592 22710
rect 5540 22646 5592 22652
rect 5736 22642 5764 23054
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 5540 21548 5592 21554
rect 5540 21490 5592 21496
rect 5552 20398 5580 21490
rect 5644 20466 5672 22374
rect 6012 21622 6040 23462
rect 6000 21616 6052 21622
rect 6000 21558 6052 21564
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5552 19446 5580 20334
rect 5540 19440 5592 19446
rect 5540 19382 5592 19388
rect 5552 18766 5580 19382
rect 5644 18834 5672 20402
rect 5828 19854 5856 20946
rect 6104 20942 6132 23666
rect 6196 22681 6224 24074
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6182 22672 6238 22681
rect 6182 22607 6238 22616
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 21010 6224 22442
rect 6288 21146 6316 23666
rect 6380 23662 6408 25230
rect 6472 25226 6500 26182
rect 6656 25906 6684 26318
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6748 26042 6776 26182
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6552 25764 6604 25770
rect 6552 25706 6604 25712
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6366 22672 6422 22681
rect 6366 22607 6368 22616
rect 6420 22607 6422 22616
rect 6368 22578 6420 22584
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 6092 20936 6144 20942
rect 6090 20904 6092 20913
rect 6144 20904 6146 20913
rect 6380 20874 6408 22578
rect 6472 21554 6500 25162
rect 6564 23730 6592 25706
rect 6748 25378 6776 25978
rect 6932 25906 6960 26726
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 7012 25764 7064 25770
rect 7012 25706 7064 25712
rect 6656 25350 6776 25378
rect 6656 24818 6684 25350
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6748 24834 6776 25230
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 6840 24954 6868 25094
rect 6828 24948 6880 24954
rect 6828 24890 6880 24896
rect 6644 24812 6696 24818
rect 6748 24806 6868 24834
rect 6644 24754 6696 24760
rect 6736 24336 6788 24342
rect 6736 24278 6788 24284
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6748 22710 6776 24278
rect 6840 23526 6868 24806
rect 7024 24750 7052 25706
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 7116 24954 7144 25638
rect 7208 25294 7236 26182
rect 7484 25838 7512 27406
rect 7576 27130 7604 28494
rect 8024 28416 8076 28422
rect 8024 28358 8076 28364
rect 8036 28150 8064 28358
rect 8024 28144 8076 28150
rect 8024 28086 8076 28092
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7760 27577 7788 27950
rect 7746 27568 7802 27577
rect 8220 27538 8248 28494
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 9048 28150 9076 28358
rect 9036 28144 9088 28150
rect 9036 28086 9088 28092
rect 9140 27878 9168 28494
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 7746 27503 7802 27512
rect 8208 27532 8260 27538
rect 7656 27328 7708 27334
rect 7654 27296 7656 27305
rect 7708 27296 7710 27305
rect 7654 27231 7710 27240
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 7668 26246 7696 27231
rect 7760 26994 7788 27503
rect 8208 27474 8260 27480
rect 9140 27470 9168 27814
rect 8484 27464 8536 27470
rect 7838 27432 7894 27441
rect 8484 27406 8536 27412
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 7838 27367 7840 27376
rect 7892 27367 7894 27376
rect 8024 27396 8076 27402
rect 7840 27338 7892 27344
rect 8024 27338 8076 27344
rect 8036 27062 8064 27338
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8128 27062 8156 27270
rect 8496 27130 8524 27406
rect 9128 27328 9180 27334
rect 9128 27270 9180 27276
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 9140 27062 9168 27270
rect 8024 27056 8076 27062
rect 8024 26998 8076 27004
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 9128 27056 9180 27062
rect 9128 26998 9180 27004
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 8484 26444 8536 26450
rect 8484 26386 8536 26392
rect 8496 26330 8524 26386
rect 8404 26302 8524 26330
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 7656 26240 7708 26246
rect 7656 26182 7708 26188
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8312 25974 8340 26182
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 7576 25294 7604 25842
rect 7656 25696 7708 25702
rect 7656 25638 7708 25644
rect 7668 25294 7696 25638
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7656 25288 7708 25294
rect 7656 25230 7708 25236
rect 7380 25152 7432 25158
rect 7760 25106 7788 25842
rect 7380 25094 7432 25100
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 7392 24886 7420 25094
rect 7668 25078 7788 25106
rect 7380 24880 7432 24886
rect 7380 24822 7432 24828
rect 7012 24744 7064 24750
rect 7012 24686 7064 24692
rect 7668 24682 7696 25078
rect 7852 24886 7880 25842
rect 8404 25770 8432 26302
rect 8392 25764 8444 25770
rect 8392 25706 8444 25712
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7944 25430 7972 25638
rect 7932 25424 7984 25430
rect 7932 25366 7984 25372
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 7564 24676 7616 24682
rect 7564 24618 7616 24624
rect 7656 24676 7708 24682
rect 7656 24618 7708 24624
rect 7576 24410 7604 24618
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7668 23866 7696 24618
rect 7852 24410 7880 24822
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7748 24200 7800 24206
rect 7800 24160 7880 24188
rect 7748 24142 7800 24148
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7196 23724 7248 23730
rect 7196 23666 7248 23672
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6736 22704 6788 22710
rect 6736 22646 6788 22652
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6564 22166 6592 22510
rect 6552 22160 6604 22166
rect 6552 22102 6604 22108
rect 6748 22030 6776 22646
rect 6840 22098 6868 23462
rect 7208 23254 7236 23666
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7196 23248 7248 23254
rect 7196 23190 7248 23196
rect 6920 22704 6972 22710
rect 6920 22646 6972 22652
rect 6932 22506 6960 22646
rect 6920 22500 6972 22506
rect 6920 22442 6972 22448
rect 7208 22166 7236 23190
rect 7392 23118 7420 23530
rect 7380 23112 7432 23118
rect 7472 23112 7524 23118
rect 7380 23054 7432 23060
rect 7470 23080 7472 23089
rect 7576 23100 7604 23666
rect 7524 23080 7604 23100
rect 7526 23072 7604 23080
rect 7470 23015 7526 23024
rect 7656 23044 7708 23050
rect 7708 23004 7788 23032
rect 7656 22986 7708 22992
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7380 22432 7432 22438
rect 7380 22374 7432 22380
rect 7196 22160 7248 22166
rect 7196 22102 7248 22108
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 6736 22024 6788 22030
rect 6736 21966 6788 21972
rect 6828 21956 6880 21962
rect 6880 21916 6960 21944
rect 6828 21898 6880 21904
rect 6552 21888 6604 21894
rect 6550 21856 6552 21865
rect 6604 21856 6606 21865
rect 6550 21791 6606 21800
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 6656 21554 6684 21626
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6656 21418 6684 21490
rect 6552 21412 6604 21418
rect 6552 21354 6604 21360
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6564 20942 6592 21354
rect 6828 21344 6880 21350
rect 6828 21286 6880 21292
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6552 20936 6604 20942
rect 6604 20896 6684 20924
rect 6552 20878 6604 20884
rect 6090 20839 6146 20848
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 6000 20800 6052 20806
rect 6000 20742 6052 20748
rect 5920 20262 5948 20742
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5736 18222 5764 18838
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5356 18148 5408 18154
rect 5356 18090 5408 18096
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5368 16114 5396 17750
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5460 15706 5488 16118
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5460 14074 5488 14282
rect 5552 14278 5580 18090
rect 5736 17746 5764 18158
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5736 17338 5764 17682
rect 6012 17678 6040 20742
rect 6196 20398 6224 20810
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6196 20058 6224 20334
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6380 19854 6408 20198
rect 6472 19990 6500 20878
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6564 19854 6592 20742
rect 6656 19922 6684 20896
rect 6748 19990 6776 21082
rect 6840 20942 6868 21286
rect 6932 21026 6960 21916
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 6932 21010 7052 21026
rect 6920 21004 7052 21010
rect 6972 20998 7052 21004
rect 6920 20946 6972 20952
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20602 6868 20878
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6932 20466 6960 20810
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 7024 19802 7052 20998
rect 7116 20534 7144 21830
rect 7208 21486 7236 22102
rect 7392 22030 7420 22374
rect 7668 22098 7696 22646
rect 7760 22642 7788 23004
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7760 22506 7788 22578
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7656 22092 7708 22098
rect 7656 22034 7708 22040
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7288 21956 7340 21962
rect 7288 21898 7340 21904
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7300 20942 7328 21898
rect 7392 21350 7420 21966
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7484 21146 7512 22034
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 6288 18698 6316 19790
rect 6460 19780 6512 19786
rect 7024 19774 7144 19802
rect 6460 19722 6512 19728
rect 6472 18970 6500 19722
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 7024 19378 7052 19654
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7012 19372 7064 19378
rect 7012 19314 7064 19320
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6748 18698 6776 19314
rect 6932 18970 6960 19314
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6288 17882 6316 18634
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5736 16726 5764 17274
rect 5724 16720 5776 16726
rect 5724 16662 5776 16668
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5644 15434 5672 15982
rect 5736 15978 5764 16662
rect 6012 16250 6040 17614
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 17338 6960 17546
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6840 16658 6868 17138
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 7024 16522 7052 19178
rect 7116 18766 7144 19774
rect 7208 18970 7236 20334
rect 7484 20074 7512 21082
rect 7392 20046 7512 20074
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7300 18970 7328 19790
rect 7392 19378 7420 20046
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19514 7512 19858
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7380 19372 7432 19378
rect 7668 19334 7696 22034
rect 7746 21856 7802 21865
rect 7852 21842 7880 24160
rect 7944 24138 7972 25366
rect 8404 25362 8432 25706
rect 8392 25356 8444 25362
rect 8392 25298 8444 25304
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7944 22420 7972 24074
rect 8036 23866 8064 25162
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 8128 24206 8156 25094
rect 8208 24404 8260 24410
rect 8208 24346 8260 24352
rect 8220 24274 8248 24346
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8116 24200 8168 24206
rect 8116 24142 8168 24148
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 8036 23730 8064 23802
rect 8588 23730 8616 26318
rect 9232 25906 9260 29582
rect 9312 28756 9364 28762
rect 9312 28698 9364 28704
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9232 25498 9260 25842
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8680 24886 8708 25230
rect 8668 24880 8720 24886
rect 8668 24822 8720 24828
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8680 24206 8708 24686
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8760 24336 8812 24342
rect 8760 24278 8812 24284
rect 8668 24200 8720 24206
rect 8668 24142 8720 24148
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8668 23724 8720 23730
rect 8668 23666 8720 23672
rect 8312 23594 8616 23610
rect 8300 23588 8628 23594
rect 8352 23582 8576 23588
rect 8300 23530 8352 23536
rect 8576 23530 8628 23536
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 8036 22778 8064 23054
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 7944 22392 8064 22420
rect 7802 21814 7880 21842
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7746 21791 7802 21800
rect 7380 19314 7432 19320
rect 7576 19306 7696 19334
rect 7760 19310 7788 21791
rect 7944 21690 7972 21830
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 19922 7880 20198
rect 7944 20058 7972 20266
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7944 19802 7972 19994
rect 8036 19938 8064 22392
rect 8128 20466 8156 22578
rect 8220 22574 8248 22714
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8220 22098 8248 22510
rect 8680 22098 8708 23666
rect 8208 22092 8260 22098
rect 8208 22034 8260 22040
rect 8484 22092 8536 22098
rect 8484 22034 8536 22040
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8300 22024 8352 22030
rect 8220 21972 8300 21978
rect 8220 21966 8352 21972
rect 8220 21950 8340 21966
rect 8392 21956 8444 21962
rect 8220 21010 8248 21950
rect 8392 21898 8444 21904
rect 8404 21690 8432 21898
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8404 21554 8432 21626
rect 8496 21622 8524 22034
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8128 20330 8156 20402
rect 8404 20330 8432 20878
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8392 20324 8444 20330
rect 8392 20266 8444 20272
rect 8036 19910 8248 19938
rect 8496 19922 8524 21558
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8588 20534 8616 21490
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8680 21146 8708 21286
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8220 19854 8248 19910
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 7852 19774 7972 19802
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17338 7144 17478
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7300 16590 7328 18702
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6012 16114 6040 16186
rect 6656 16182 6684 16390
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 6644 16040 6696 16046
rect 6644 15982 6696 15988
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 6656 15706 6684 15982
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 7300 15434 7328 16526
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5552 14006 5580 14214
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 12374 5488 13874
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5552 12442 5580 12854
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5644 11898 5672 15370
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6012 13938 6040 14350
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 14074 6224 14214
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 6012 12442 6040 12718
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6104 12238 6132 13126
rect 6288 12918 6316 13194
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6288 12238 6316 12854
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6380 12170 6408 14282
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6564 12850 6592 13194
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6564 12306 6592 12786
rect 6656 12442 6684 14962
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6748 14618 6776 14758
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 14414 6868 14554
rect 6932 14550 6960 14758
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6932 14006 6960 14486
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6840 12986 6868 13874
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12889 6868 12922
rect 6826 12880 6882 12889
rect 6736 12844 6788 12850
rect 6826 12815 6882 12824
rect 6736 12786 6788 12792
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5368 10470 5396 11562
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11218 6316 11494
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6288 11082 6316 11154
rect 6748 11150 6776 12786
rect 7024 12782 7052 14010
rect 7116 13734 7144 14962
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7208 13326 7236 13806
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12850 7236 13262
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7300 12850 7328 13194
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 11620 7248 11626
rect 7196 11562 7248 11568
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 6656 10742 6684 10950
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 7116 10674 7144 10950
rect 7208 10810 7236 11562
rect 7300 10826 7328 12378
rect 7392 11014 7420 14418
rect 7484 12442 7512 18702
rect 7576 17678 7604 19306
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7576 17338 7604 17614
rect 7852 17610 7880 19774
rect 7932 19712 7984 19718
rect 7930 19680 7932 19689
rect 8024 19712 8076 19718
rect 7984 19680 7986 19689
rect 8024 19654 8076 19660
rect 7930 19615 7986 19624
rect 8036 19446 8064 19654
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 8128 19334 8156 19790
rect 8036 19306 8156 19334
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7668 17134 7696 17274
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7668 15570 7696 17070
rect 7852 17066 7880 17546
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 12850 7604 13126
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7668 12730 7696 13262
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7576 12702 7696 12730
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7576 12322 7604 12702
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12442 7696 12582
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7484 12294 7604 12322
rect 7484 11898 7512 12294
rect 7760 12238 7788 13126
rect 7852 12986 7880 15030
rect 7932 13320 7984 13326
rect 7932 13262 7984 13268
rect 7944 12986 7972 13262
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 7852 12186 7880 12582
rect 7944 12306 7972 12786
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7576 11762 7604 12174
rect 7852 12158 7972 12186
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11830 7880 12038
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11354 7604 11698
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7196 10804 7248 10810
rect 7300 10798 7420 10826
rect 7196 10746 7248 10752
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5368 10198 5396 10406
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5460 10062 5488 10406
rect 5736 10266 5764 10542
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5276 9646 5396 9674
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2700 8974 2728 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9042 4660 9318
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2976 7342 3004 7822
rect 3160 7342 3188 8978
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8514 5396 9646
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6012 8906 6040 9590
rect 6380 9042 6408 10066
rect 6564 10062 6592 10610
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5276 8486 5396 8514
rect 5632 8492 5684 8498
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2976 7002 3004 7278
rect 2964 6996 3016 7002
rect 2964 6938 3016 6944
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2424 6458 2452 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1950 5808 2006 5817
rect 3160 5778 3188 7278
rect 4448 7274 4476 7754
rect 4436 7268 4488 7274
rect 4436 7210 4488 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6866 4660 7142
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 1950 5743 2006 5752
rect 3148 5772 3200 5778
rect 3148 5714 3200 5720
rect 4080 5692 4108 6802
rect 4724 6798 4752 7958
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7528 4844 7890
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4816 7500 4936 7528
rect 4908 7410 4936 7500
rect 5276 7449 5304 8486
rect 5632 8434 5684 8440
rect 5262 7440 5318 7449
rect 4896 7404 4948 7410
rect 5262 7375 5318 7384
rect 4896 7346 4948 7352
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5704 4212 5710
rect 4080 5664 4160 5692
rect 4160 5646 4212 5652
rect 4172 5234 4200 5646
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4448 5370 4476 5578
rect 4816 5370 4844 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4436 5364 4488 5370
rect 4436 5306 4488 5312
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 5460 5166 5488 5714
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5552 5370 5580 5646
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5644 5234 5672 8434
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5908 7948 5960 7954
rect 5960 7908 6132 7936
rect 5908 7890 5960 7896
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5736 7410 5764 7822
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5828 7324 5856 7890
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5828 7296 5948 7324
rect 5920 7154 5948 7296
rect 6012 7274 6040 7686
rect 6104 7478 6132 7908
rect 6380 7818 6408 8978
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6196 7154 6224 7346
rect 5920 7126 6224 7154
rect 5920 5574 5948 7126
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5920 5302 5948 5510
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5644 5098 5672 5170
rect 6368 5160 6420 5166
rect 6472 5148 6500 8774
rect 6564 7546 6592 9998
rect 7024 9674 7052 10202
rect 6932 9646 7052 9674
rect 6932 9586 6960 9646
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6644 9376 6696 9382
rect 6642 9344 6644 9353
rect 6696 9344 6698 9353
rect 6642 9279 6698 9288
rect 6748 9178 6776 9522
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 8430 6868 9386
rect 7024 9382 7052 9646
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6932 8498 6960 9318
rect 7116 8906 7144 10610
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7208 9994 7236 10474
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7208 9654 7236 9930
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8634 7236 8842
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 7886 6868 8366
rect 7300 8090 7328 9862
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 7288 7880 7340 7886
rect 7392 7857 7420 10798
rect 7668 10266 7696 11630
rect 7760 10810 7788 11630
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7944 10470 7972 12158
rect 8036 11626 8064 19306
rect 8220 18834 8248 19790
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8312 18630 8340 19722
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8404 18766 8432 19314
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8312 17202 8340 17818
rect 8496 17678 8524 19858
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8404 17134 8432 17478
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16726 8432 17070
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 16182 8248 16526
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 15502 8524 15846
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 13938 8340 14894
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12238 8156 13262
rect 8220 12850 8248 13738
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8024 11620 8076 11626
rect 8024 11562 8076 11568
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10266 7972 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7470 9344 7526 9353
rect 7470 9279 7526 9288
rect 7484 8430 7512 9279
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8566 7604 9114
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7288 7822 7340 7828
rect 7378 7848 7434 7857
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7342 6684 7686
rect 7116 7410 7144 7686
rect 7300 7478 7328 7822
rect 7378 7783 7434 7792
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6564 6322 6592 7210
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6656 6254 6684 7278
rect 6840 6934 6868 7346
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 7024 5710 7052 6122
rect 7392 5710 7420 7346
rect 7484 5778 7512 8366
rect 7576 7818 7604 8502
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 7002 7788 7142
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7852 6866 7880 9998
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 7886 8064 8230
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7410 7972 7686
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6656 5302 6684 5510
rect 8036 5370 8064 5646
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6420 5120 6500 5148
rect 6368 5102 6420 5108
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 6380 4146 6408 5102
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 8128 2774 8156 12174
rect 8220 11558 8248 12650
rect 8312 12238 8340 13874
rect 8496 13258 8524 14418
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 12889 8524 13194
rect 8482 12880 8538 12889
rect 8482 12815 8484 12824
rect 8536 12815 8538 12824
rect 8484 12786 8536 12792
rect 8588 12434 8616 20470
rect 8772 19802 8800 24278
rect 8852 24268 8904 24274
rect 8852 24210 8904 24216
rect 8680 19774 8800 19802
rect 8680 19514 8708 19774
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8772 19514 8800 19654
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8680 19174 8708 19314
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18902 8708 19110
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8864 17218 8892 24210
rect 8956 24206 8984 24550
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 8956 20874 8984 22578
rect 9232 22094 9260 25434
rect 9324 23186 9352 28698
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9416 25770 9444 26318
rect 9404 25764 9456 25770
rect 9404 25706 9456 25712
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9312 23180 9364 23186
rect 9312 23122 9364 23128
rect 9048 22066 9260 22094
rect 9312 22094 9364 22098
rect 9416 22094 9444 23666
rect 9312 22092 9444 22094
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8956 20058 8984 20402
rect 9048 20330 9076 22066
rect 9364 22066 9444 22092
rect 9312 22034 9364 22040
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9140 21418 9168 21966
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9324 21146 9352 22034
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9416 21554 9444 21898
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9232 20466 9260 20878
rect 9324 20602 9352 20878
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9036 20324 9088 20330
rect 9036 20266 9088 20272
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9140 19786 9168 20402
rect 9232 20369 9260 20402
rect 9416 20398 9444 21490
rect 9508 21434 9536 30058
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 10416 28620 10468 28626
rect 10416 28562 10468 28568
rect 10428 28506 10456 28562
rect 10244 28478 10456 28506
rect 11164 28490 11192 28970
rect 10508 28484 10560 28490
rect 10244 28082 10272 28478
rect 10508 28426 10560 28432
rect 11152 28484 11204 28490
rect 11152 28426 11204 28432
rect 10520 28218 10548 28426
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10692 28212 10744 28218
rect 10692 28154 10744 28160
rect 10048 28076 10100 28082
rect 10048 28018 10100 28024
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10060 27674 10088 28018
rect 10048 27668 10100 27674
rect 10048 27610 10100 27616
rect 10152 27538 10180 28018
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 10244 27470 10272 28018
rect 10704 27606 10732 28154
rect 11348 28082 11376 28358
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10796 27674 10824 27814
rect 10784 27668 10836 27674
rect 10784 27610 10836 27616
rect 10692 27600 10744 27606
rect 10692 27542 10744 27548
rect 10048 27464 10100 27470
rect 10048 27406 10100 27412
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 9586 27296 9642 27305
rect 9586 27231 9642 27240
rect 9600 27130 9628 27231
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 10060 26790 10088 27406
rect 11072 27402 11100 27882
rect 10968 27396 11020 27402
rect 10968 27338 11020 27344
rect 11060 27396 11112 27402
rect 11060 27338 11112 27344
rect 10980 26994 11008 27338
rect 10968 26988 11020 26994
rect 10968 26930 11020 26936
rect 11164 26926 11192 28018
rect 11348 27470 11376 28018
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9864 26240 9916 26246
rect 9864 26182 9916 26188
rect 9876 25906 9904 26182
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9692 25294 9720 25434
rect 9784 25294 9812 25774
rect 9864 25764 9916 25770
rect 9864 25706 9916 25712
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9600 23730 9628 24822
rect 9784 24206 9812 25094
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9770 23760 9826 23769
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9680 23724 9732 23730
rect 9770 23695 9772 23704
rect 9680 23666 9732 23672
rect 9824 23695 9826 23704
rect 9772 23666 9824 23672
rect 9692 22778 9720 23666
rect 9772 23520 9824 23526
rect 9772 23462 9824 23468
rect 9784 23254 9812 23462
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9600 21554 9628 21830
rect 9784 21729 9812 22034
rect 9770 21720 9826 21729
rect 9770 21655 9826 21664
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9508 21406 9628 21434
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 9508 20602 9536 20878
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9404 20392 9456 20398
rect 9218 20360 9274 20369
rect 9404 20334 9456 20340
rect 9218 20295 9274 20304
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9508 19922 9536 20266
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9128 19440 9180 19446
rect 9128 19382 9180 19388
rect 9402 19408 9458 19417
rect 9140 19174 9168 19382
rect 9402 19343 9404 19352
rect 9456 19343 9458 19352
rect 9404 19314 9456 19320
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 8944 18760 8996 18766
rect 8944 18702 8996 18708
rect 8956 18154 8984 18702
rect 9140 18698 9168 19110
rect 9128 18692 9180 18698
rect 9128 18634 9180 18640
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8956 17882 8984 18090
rect 9140 17921 9168 18634
rect 9126 17912 9182 17921
rect 8944 17876 8996 17882
rect 9126 17847 9182 17856
rect 8944 17818 8996 17824
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8772 17190 8892 17218
rect 8772 12442 8800 17190
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8864 16114 8892 16594
rect 9140 16250 9168 17478
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8956 15706 8984 15982
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9048 15502 9076 16118
rect 9140 15502 9168 16186
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 9140 13938 9168 14826
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9232 13938 9260 14418
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 12850 9076 13670
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8760 12436 8812 12442
rect 8588 12406 8708 12434
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11898 8340 12038
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8220 7546 8248 7822
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7546 8340 7686
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8220 6458 8248 7346
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 6866 8432 7142
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8496 6798 8524 7754
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8588 7002 8616 7346
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8312 5914 8340 6734
rect 8496 6458 8524 6734
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8588 5846 8616 6258
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8496 5370 8524 5646
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8588 5302 8616 5782
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8036 2746 8156 2774
rect 4988 2576 5040 2582
rect 4986 2544 4988 2553
rect 5040 2544 5042 2553
rect 4986 2479 5042 2488
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 952 2145 980 2382
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 938 2136 994 2145
rect 938 2071 994 2080
rect 1596 1970 1624 2246
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 846 912 902 921
rect 846 847 902 856
rect 1964 800 1992 2382
rect 3252 800 3280 2382
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4540 800 4568 2314
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5828 800 5856 2382
rect 7116 800 7144 2382
rect 7760 800 7788 2382
rect 8036 2310 8064 2746
rect 8680 2650 8708 12406
rect 8760 12378 8812 12384
rect 8864 11830 8892 12786
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12646 8984 12718
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12170 8984 12582
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8864 11150 8892 11766
rect 8956 11626 8984 12106
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9048 11762 9076 12038
rect 9416 11880 9444 19314
rect 9508 18970 9536 19722
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9508 18766 9536 18906
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9508 12850 9536 13126
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9600 12434 9628 21406
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20534 9720 20810
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9692 19786 9720 20470
rect 9876 20398 9904 25706
rect 9956 25696 10008 25702
rect 9956 25638 10008 25644
rect 9968 25498 9996 25638
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 10060 24818 10088 26726
rect 10336 26382 10364 26862
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10324 26376 10376 26382
rect 11244 26376 11296 26382
rect 10376 26324 10640 26330
rect 10324 26318 10640 26324
rect 11244 26318 11296 26324
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9968 24410 9996 24550
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9968 24206 9996 24346
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 9968 23526 9996 24006
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 10060 23118 10088 24006
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9968 22030 9996 22714
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 9968 21146 9996 21422
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9956 20936 10008 20942
rect 10060 20924 10088 23054
rect 10008 20896 10088 20924
rect 9956 20878 10008 20884
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 9864 20392 9916 20398
rect 9864 20334 9916 20340
rect 9784 19854 9812 20334
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9680 19780 9732 19786
rect 9680 19722 9732 19728
rect 9876 19446 9904 19994
rect 9864 19440 9916 19446
rect 9784 19388 9864 19394
rect 9784 19382 9916 19388
rect 9784 19366 9904 19382
rect 9680 18896 9732 18902
rect 9678 18864 9680 18873
rect 9732 18864 9734 18873
rect 9678 18799 9734 18808
rect 9692 18698 9720 18799
rect 9784 18766 9812 19366
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 18766 9904 19246
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9876 18578 9904 18702
rect 9784 18550 9904 18578
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 16114 9720 17138
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9784 15994 9812 18550
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9876 16590 9904 17546
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9692 15966 9812 15994
rect 9692 15162 9720 15966
rect 9876 15910 9904 16526
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9784 15570 9812 15846
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9876 15434 9904 15846
rect 9864 15428 9916 15434
rect 9864 15370 9916 15376
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9784 12968 9812 15302
rect 9784 12940 9904 12968
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9232 11852 9444 11880
rect 9508 12406 9628 12434
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 9140 11354 9168 11698
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8864 10470 8892 10678
rect 8956 10674 8984 10746
rect 9140 10674 9168 10950
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8772 10062 8800 10406
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 9048 9722 9076 10610
rect 9232 9738 9260 11852
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9324 11626 9352 11698
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9324 11150 9352 11290
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9416 10674 9444 11698
rect 9508 11540 9536 12406
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9600 11608 9628 12242
rect 9680 12232 9732 12238
rect 9678 12200 9680 12209
rect 9732 12200 9734 12209
rect 9678 12135 9734 12144
rect 9784 11898 9812 12786
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11694 9904 12940
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9680 11620 9732 11626
rect 9600 11580 9680 11608
rect 9680 11562 9732 11568
rect 9508 11512 9628 11540
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9508 11150 9536 11222
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9324 10470 9352 10610
rect 9508 10606 9536 11086
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9140 9710 9260 9738
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8864 9042 8892 9454
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5778 8800 6122
rect 8760 5772 8812 5778
rect 8760 5714 8812 5720
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8864 4826 8892 5578
rect 8956 5234 8984 5646
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8220 2530 8248 2586
rect 8220 2514 8340 2530
rect 8220 2508 8352 2514
rect 8220 2502 8300 2508
rect 8300 2450 8352 2456
rect 8864 2446 8892 4762
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8956 2378 8984 5170
rect 9048 5098 9076 8978
rect 9140 8634 9168 9710
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 8974 9260 9522
rect 9416 8974 9444 9590
rect 9508 9518 9536 10542
rect 9600 9518 9628 11512
rect 9692 11206 9904 11234
rect 9692 11082 9720 11206
rect 9876 11150 9904 11206
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10674 9720 11018
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10810 9812 10950
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9968 10554 9996 20878
rect 10048 20528 10100 20534
rect 10048 20470 10100 20476
rect 10060 19854 10088 20470
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 18578 10088 19790
rect 10152 18698 10180 26318
rect 10336 26314 10640 26318
rect 10336 26308 10652 26314
rect 10336 26302 10600 26308
rect 10600 26250 10652 26256
rect 10876 26308 10928 26314
rect 10876 26250 10928 26256
rect 10888 26042 10916 26250
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10980 25906 11008 26182
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 10692 25832 10744 25838
rect 10692 25774 10744 25780
rect 10704 25430 10732 25774
rect 10692 25424 10744 25430
rect 10692 25366 10744 25372
rect 11256 25362 11284 26318
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10232 24676 10284 24682
rect 10232 24618 10284 24624
rect 10244 24274 10272 24618
rect 10428 24274 10456 25162
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10232 24268 10284 24274
rect 10416 24268 10468 24274
rect 10284 24228 10364 24256
rect 10232 24210 10284 24216
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10244 23594 10272 24006
rect 10232 23588 10284 23594
rect 10232 23530 10284 23536
rect 10244 23118 10272 23530
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10336 22642 10364 24228
rect 10416 24210 10468 24216
rect 10520 24138 10548 24754
rect 10612 24138 10640 25230
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10600 24132 10652 24138
rect 10600 24074 10652 24080
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10336 22409 10364 22578
rect 10520 22574 10548 24074
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10322 22400 10378 22409
rect 10322 22335 10378 22344
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10244 21690 10272 22102
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10336 21894 10364 21966
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10520 21350 10548 22034
rect 10612 22030 10640 23190
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10612 21554 10640 21626
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10704 20534 10732 25230
rect 11164 24614 11192 25230
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10796 23730 10824 24006
rect 11152 23792 11204 23798
rect 11150 23760 11152 23769
rect 11204 23760 11206 23769
rect 10784 23724 10836 23730
rect 11150 23695 11206 23704
rect 10784 23666 10836 23672
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10888 22778 10916 23122
rect 11072 23118 11100 23462
rect 11164 23118 11192 23695
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 11256 23322 11284 23462
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11256 23118 11284 23258
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10796 20602 10824 22374
rect 10888 22012 10916 22578
rect 10968 22024 11020 22030
rect 10888 21984 10968 22012
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10244 19310 10272 20402
rect 10796 19854 10824 20538
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 10612 19514 10640 19722
rect 10704 19514 10732 19790
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10520 18970 10548 19314
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10324 18624 10376 18630
rect 10060 18550 10180 18578
rect 10324 18566 10376 18572
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16114 10088 16390
rect 10152 16130 10180 18550
rect 10336 18222 10364 18566
rect 10428 18358 10456 18702
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10888 18222 10916 21984
rect 10968 21966 11020 21972
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11256 21894 11284 21966
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21418 11284 21830
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 11348 20874 11376 27406
rect 11624 24138 11652 30126
rect 12072 30116 12124 30122
rect 12072 30058 12124 30064
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 11716 22438 11744 26386
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11900 25498 11928 25842
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11992 24206 12020 24550
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11704 22432 11756 22438
rect 11426 22400 11482 22409
rect 11704 22374 11756 22380
rect 11426 22335 11482 22344
rect 11440 21962 11468 22335
rect 11716 22166 11744 22374
rect 11704 22160 11756 22166
rect 11704 22102 11756 22108
rect 12084 22094 12112 30058
rect 12164 30048 12216 30054
rect 12164 29990 12216 29996
rect 12532 30048 12584 30054
rect 12532 29990 12584 29996
rect 13544 30048 13596 30054
rect 13544 29990 13596 29996
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 15660 30048 15712 30054
rect 15660 29990 15712 29996
rect 12176 24206 12204 29990
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12348 28552 12400 28558
rect 12348 28494 12400 28500
rect 12360 27946 12388 28494
rect 12348 27940 12400 27946
rect 12348 27882 12400 27888
rect 12452 26994 12480 29106
rect 12544 29073 12572 29990
rect 13556 29646 13584 29990
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13084 29504 13136 29510
rect 13084 29446 13136 29452
rect 12624 29096 12676 29102
rect 12530 29064 12586 29073
rect 12624 29038 12676 29044
rect 12530 28999 12586 29008
rect 12636 28082 12664 29038
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12728 28218 12756 28494
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12912 28150 12940 28358
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12624 27396 12676 27402
rect 12624 27338 12676 27344
rect 12636 27130 12664 27338
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12624 26852 12676 26858
rect 12624 26794 12676 26800
rect 12636 26518 12664 26794
rect 12624 26512 12676 26518
rect 12624 26454 12676 26460
rect 13096 26382 13124 29446
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13648 28558 13676 29106
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13188 28218 13216 28494
rect 14004 28484 14056 28490
rect 14004 28426 14056 28432
rect 13636 28416 13688 28422
rect 13636 28358 13688 28364
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13188 27606 13216 28154
rect 13648 28150 13676 28358
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13636 28144 13688 28150
rect 13636 28086 13688 28092
rect 13176 27600 13228 27606
rect 13176 27542 13228 27548
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13280 26994 13308 27270
rect 13268 26988 13320 26994
rect 13268 26930 13320 26936
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 26450 13216 26726
rect 13176 26444 13228 26450
rect 13176 26386 13228 26392
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12452 26042 12480 26182
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12268 25430 12296 25842
rect 12728 25786 12756 26182
rect 12912 25906 12940 26318
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 12636 25758 12756 25786
rect 12808 25764 12860 25770
rect 12636 25702 12664 25758
rect 12808 25706 12860 25712
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12256 24744 12308 24750
rect 12256 24686 12308 24692
rect 12268 24206 12296 24686
rect 12164 24200 12216 24206
rect 12256 24200 12308 24206
rect 12164 24142 12216 24148
rect 12254 24168 12256 24177
rect 12308 24168 12310 24177
rect 12176 22574 12204 24142
rect 12254 24103 12310 24112
rect 12256 23316 12308 23322
rect 12256 23258 12308 23264
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 11992 22066 12112 22094
rect 11612 22024 11664 22030
rect 11664 21972 11744 21978
rect 11612 21966 11744 21972
rect 11428 21956 11480 21962
rect 11624 21950 11744 21966
rect 11992 21962 12020 22066
rect 12072 22024 12124 22030
rect 12176 22012 12204 22510
rect 12124 21984 12204 22012
rect 12072 21966 12124 21972
rect 11428 21898 11480 21904
rect 11716 21894 11744 21950
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11532 21078 11560 21830
rect 11624 21690 11652 21830
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11612 21548 11664 21554
rect 11612 21490 11664 21496
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 10980 20466 11008 20810
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11336 20460 11388 20466
rect 11336 20402 11388 20408
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11256 19854 11284 19994
rect 11348 19990 11376 20402
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11532 20058 11560 20198
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11336 19984 11388 19990
rect 11336 19926 11388 19932
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10980 18902 11008 19314
rect 11532 19310 11560 19994
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10230 17504 10286 17513
rect 10230 17439 10286 17448
rect 10244 17338 10272 17439
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10244 16232 10272 17138
rect 10336 16658 10364 18158
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10428 17338 10456 18022
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10428 17202 10456 17274
rect 10704 17202 10732 17818
rect 10796 17678 10824 18022
rect 10980 17678 11008 18226
rect 11072 17746 11100 18362
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10612 17082 10640 17138
rect 10796 17082 10824 17478
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10980 17202 11008 17274
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 10612 17054 10824 17082
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10324 16244 10376 16250
rect 10244 16204 10324 16232
rect 10324 16186 10376 16192
rect 10048 16108 10100 16114
rect 10152 16102 10732 16130
rect 10796 16114 10824 17054
rect 10980 16590 11008 17138
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16114 11008 16390
rect 10048 16050 10100 16056
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10060 15706 10088 15914
rect 10336 15858 10364 15914
rect 10244 15830 10364 15858
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10244 15502 10272 15830
rect 10520 15706 10548 15982
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10336 15502 10364 15642
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10152 15026 10180 15098
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10060 14414 10088 14486
rect 10152 14414 10180 14758
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10336 14074 10364 14486
rect 10612 14414 10640 14486
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 12986 10364 14010
rect 10520 13938 10548 14214
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10244 12714 10272 12854
rect 10336 12850 10364 12922
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10428 12782 10456 13738
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10232 12708 10284 12714
rect 10232 12650 10284 12656
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10060 12442 10088 12582
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10152 12238 10180 12582
rect 10244 12238 10272 12650
rect 10520 12442 10548 13670
rect 10612 13326 10640 14214
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10508 12436 10560 12442
rect 10704 12434 10732 16102
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10980 15706 11008 16050
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11348 15502 11376 17138
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11624 15162 11652 21490
rect 11900 21434 11928 21898
rect 11992 21554 12020 21898
rect 12070 21720 12126 21729
rect 12070 21655 12126 21664
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11716 21406 11928 21434
rect 11716 20641 11744 21406
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20942 11928 21286
rect 11888 20936 11940 20942
rect 11888 20878 11940 20884
rect 11796 20868 11848 20874
rect 11796 20810 11848 20816
rect 11702 20632 11758 20641
rect 11702 20567 11758 20576
rect 11716 20534 11744 20567
rect 11704 20528 11756 20534
rect 11704 20470 11756 20476
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11716 19922 11744 20198
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11808 18290 11836 20810
rect 11888 20800 11940 20806
rect 11888 20742 11940 20748
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 16250 11744 17478
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11808 16182 11836 18226
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11808 15706 11836 15846
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 13938 10824 14418
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 12714 10824 13874
rect 10888 13326 10916 14214
rect 11072 13938 11100 14350
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10980 13802 11008 13874
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 11164 13716 11192 14962
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 11256 14006 11284 14486
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11244 14000 11296 14006
rect 11296 13960 11468 13988
rect 11244 13942 11296 13948
rect 11072 13688 11192 13716
rect 11244 13728 11296 13734
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 11072 12442 11100 13688
rect 11244 13670 11296 13676
rect 11256 13394 11284 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12436 11112 12442
rect 10704 12406 10824 12434
rect 10508 12378 10560 12384
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10152 11830 10180 12174
rect 10520 11898 10548 12174
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 11898 10732 12106
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 9968 10526 10364 10554
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10062 10272 10406
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9680 9512 9732 9518
rect 9732 9472 9812 9500
rect 9680 9454 9732 9460
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9042 9628 9318
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9416 8430 9444 8910
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9416 8022 9444 8366
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9140 6780 9168 7278
rect 9220 6792 9272 6798
rect 9140 6752 9220 6780
rect 9220 6734 9272 6740
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9140 6254 9168 6394
rect 9508 6322 9536 7822
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5098 9168 6190
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5234 9260 5646
rect 9600 5642 9628 7414
rect 9692 7410 9720 9114
rect 9784 7410 9812 9472
rect 9876 8294 9904 9998
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9784 6934 9812 7346
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 7206 9904 7278
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9968 5370 9996 9998
rect 10060 9722 10088 9998
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 10152 9518 10180 9862
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10244 9178 10272 9386
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10336 9058 10364 10526
rect 10520 10266 10548 11698
rect 10612 11354 10640 11698
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11354 10732 11562
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10612 10062 10640 10542
rect 10704 10470 10732 11154
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10152 9030 10364 9058
rect 10046 8392 10102 8401
rect 10046 8327 10102 8336
rect 10060 7886 10088 8327
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10152 6440 10180 9030
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 7410 10272 8774
rect 10336 8090 10364 8910
rect 10520 8838 10548 8910
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10336 7886 10364 7919
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10336 6798 10364 7822
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10428 7546 10456 7754
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10428 6798 10456 7482
rect 10520 7274 10548 8774
rect 10692 7336 10744 7342
rect 10690 7304 10692 7313
rect 10744 7304 10746 7313
rect 10508 7268 10560 7274
rect 10690 7239 10746 7248
rect 10508 7210 10560 7216
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10060 6412 10180 6440
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 9048 3534 9076 5034
rect 10060 4758 10088 6412
rect 10428 6390 10456 6734
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5914 10180 6258
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 4758 10180 5510
rect 10244 5234 10272 6054
rect 10324 5704 10376 5710
rect 10322 5672 10324 5681
rect 10416 5704 10468 5710
rect 10376 5672 10378 5681
rect 10416 5646 10468 5652
rect 10322 5607 10378 5616
rect 10428 5273 10456 5646
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10414 5264 10470 5273
rect 10232 5228 10284 5234
rect 10704 5234 10732 5510
rect 10414 5199 10470 5208
rect 10692 5228 10744 5234
rect 10232 5170 10284 5176
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9968 3738 9996 4150
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9600 3058 9628 3470
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 10152 2514 10180 4694
rect 10428 2650 10456 5199
rect 10692 5170 10744 5176
rect 10796 2774 10824 12406
rect 11060 12378 11112 12384
rect 11164 12238 11192 12582
rect 11348 12442 11376 13466
rect 11440 12850 11468 13960
rect 11532 13938 11560 14282
rect 11624 14006 11652 14962
rect 11900 14890 11928 20742
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 19786 12020 20402
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 12084 18426 12112 21655
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12176 19242 12204 20470
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12072 18420 12124 18426
rect 11992 18380 12072 18408
rect 11992 17746 12020 18380
rect 12072 18362 12124 18368
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12084 17882 12112 18158
rect 12268 17898 12296 23258
rect 12360 20466 12388 25094
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12622 24168 12678 24177
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12452 23186 12480 24006
rect 12544 23798 12572 24142
rect 12622 24103 12678 24112
rect 12532 23792 12584 23798
rect 12532 23734 12584 23740
rect 12636 23662 12664 24103
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12544 22030 12572 22374
rect 12728 22234 12756 22510
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12820 22094 12848 25706
rect 13004 25498 13032 26318
rect 13096 25922 13124 26318
rect 13096 25894 13216 25922
rect 13084 25832 13136 25838
rect 13084 25774 13136 25780
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13096 25430 13124 25774
rect 13188 25702 13216 25894
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13084 25424 13136 25430
rect 13084 25366 13136 25372
rect 13280 25362 13308 26930
rect 13452 26852 13504 26858
rect 13452 26794 13504 26800
rect 13464 25906 13492 26794
rect 13556 26790 13584 27270
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 13556 25922 13584 26726
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13648 26042 13676 26182
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 13452 25900 13504 25906
rect 13556 25894 13676 25922
rect 13452 25842 13504 25848
rect 13372 25498 13400 25842
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13268 25356 13320 25362
rect 13268 25298 13320 25304
rect 13464 25294 13492 25638
rect 12900 25288 12952 25294
rect 12900 25230 12952 25236
rect 13452 25288 13504 25294
rect 13452 25230 13504 25236
rect 12912 24138 12940 25230
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13268 25220 13320 25226
rect 13268 25162 13320 25168
rect 12900 24132 12952 24138
rect 12900 24074 12952 24080
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23322 13032 24074
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 13096 23730 13124 24006
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13004 22710 13032 23258
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12912 22166 12940 22374
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 13188 22094 13216 25162
rect 13280 24206 13308 25162
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13280 23662 13308 24006
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 12728 22066 12848 22094
rect 13004 22066 13216 22094
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12452 20806 12480 21898
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12360 19310 12388 20266
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12176 17870 12296 17898
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12084 16250 12112 17546
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12084 15638 12112 16186
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 12176 14074 12204 17870
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12268 17513 12296 17546
rect 12348 17536 12400 17542
rect 12254 17504 12310 17513
rect 12348 17478 12400 17484
rect 12254 17439 12310 17448
rect 12360 16998 12388 17478
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12360 15026 12388 15098
rect 12452 15026 12480 20742
rect 12544 17814 12572 21422
rect 12636 18086 12664 21422
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12728 17218 12756 22066
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12808 20936 12860 20942
rect 12808 20878 12860 20884
rect 12820 19417 12848 20878
rect 12912 20754 12940 21830
rect 13004 21554 13032 22066
rect 13280 22030 13308 22578
rect 13360 22092 13412 22098
rect 13464 22080 13492 25230
rect 13648 25226 13676 25894
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13556 23526 13584 24074
rect 13740 24070 13768 26862
rect 13924 25906 13952 28154
rect 14016 27470 14044 28426
rect 14568 28218 14596 28902
rect 14556 28212 14608 28218
rect 14556 28154 14608 28160
rect 14832 28212 14884 28218
rect 14832 28154 14884 28160
rect 14740 28144 14792 28150
rect 14740 28086 14792 28092
rect 14188 27940 14240 27946
rect 14188 27882 14240 27888
rect 14200 27674 14228 27882
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14016 27130 14044 27406
rect 14096 27396 14148 27402
rect 14096 27338 14148 27344
rect 14004 27124 14056 27130
rect 14004 27066 14056 27072
rect 14108 26994 14136 27338
rect 14384 27334 14412 27406
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14372 27328 14424 27334
rect 14372 27270 14424 27276
rect 14096 26988 14148 26994
rect 14096 26930 14148 26936
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 13924 24410 13952 25842
rect 14200 25226 14228 27270
rect 14660 26450 14688 27814
rect 14752 27674 14780 28086
rect 14740 27668 14792 27674
rect 14740 27610 14792 27616
rect 14844 27470 14872 28154
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14648 26444 14700 26450
rect 14648 26386 14700 26392
rect 14844 26042 14872 26930
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14292 25294 14320 25774
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25498 14504 25638
rect 14464 25492 14516 25498
rect 14464 25434 14516 25440
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 14188 25220 14240 25226
rect 14188 25162 14240 25168
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 13924 24274 13952 24346
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14004 24132 14056 24138
rect 14004 24074 14056 24080
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13912 23724 13964 23730
rect 13912 23666 13964 23672
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13556 22506 13584 23462
rect 13924 23254 13952 23666
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13728 22568 13780 22574
rect 13728 22510 13780 22516
rect 13544 22500 13596 22506
rect 13544 22442 13596 22448
rect 13556 22166 13584 22442
rect 13544 22160 13596 22166
rect 13544 22102 13596 22108
rect 13412 22052 13492 22080
rect 13360 22034 13412 22040
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13268 22024 13320 22030
rect 13268 21966 13320 21972
rect 13188 21729 13216 21966
rect 13174 21720 13230 21729
rect 13174 21655 13230 21664
rect 13280 21554 13308 21966
rect 13464 21622 13492 22052
rect 13740 22030 13768 22510
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13452 21616 13504 21622
rect 13452 21558 13504 21564
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13004 21146 13032 21490
rect 13280 21418 13308 21490
rect 13740 21486 13768 21966
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12912 20726 13032 20754
rect 13004 20448 13032 20726
rect 13372 20466 13400 21286
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20466 13584 20742
rect 13818 20632 13874 20641
rect 13818 20567 13874 20576
rect 13832 20534 13860 20567
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13924 20466 13952 21830
rect 13084 20460 13136 20466
rect 13004 20420 13084 20448
rect 13004 19718 13032 20420
rect 13084 20402 13136 20408
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13372 19854 13400 20402
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 12806 19408 12862 19417
rect 13188 19378 13216 19654
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 12806 19343 12862 19352
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 12544 17190 12756 17218
rect 12820 17202 12848 17546
rect 12808 17196 12860 17202
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14890 12480 14962
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11624 13734 11652 13942
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11808 13530 11836 13806
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 12452 13462 12480 13806
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11532 12442 11560 12650
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 10888 11370 10916 12174
rect 10966 11792 11022 11801
rect 10966 11727 10968 11736
rect 11020 11727 11022 11736
rect 10968 11698 11020 11704
rect 10888 11342 11008 11370
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10888 10674 10916 11222
rect 10980 11218 11008 11342
rect 11164 11286 11192 12174
rect 11256 11626 11284 12378
rect 11336 12164 11388 12170
rect 11336 12106 11388 12112
rect 11244 11620 11296 11626
rect 11244 11562 11296 11568
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11348 11082 11376 12106
rect 11624 11354 11652 13194
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11716 11762 11744 12242
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11348 10742 11376 11018
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10888 10266 10916 10610
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10980 10062 11008 10542
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9722 11008 9998
rect 11348 9994 11376 10678
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11256 8566 11284 8842
rect 11244 8560 11296 8566
rect 11244 8502 11296 8508
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8022 11008 8230
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11150 7984 11206 7993
rect 10876 7880 10928 7886
rect 11072 7834 11100 7958
rect 11150 7919 11206 7928
rect 11164 7886 11192 7919
rect 10876 7822 10928 7828
rect 10888 7478 10916 7822
rect 10980 7806 11100 7834
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10876 7472 10928 7478
rect 10876 7414 10928 7420
rect 10980 7206 11008 7806
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7410 11100 7686
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6798 11008 7142
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11072 6254 11100 7346
rect 11164 6322 11192 7822
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 10980 6100 11008 6190
rect 11256 6100 11284 7346
rect 10980 6072 11284 6100
rect 11150 5944 11206 5953
rect 11150 5879 11152 5888
rect 11204 5879 11206 5888
rect 11152 5850 11204 5856
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10968 5704 11020 5710
rect 10966 5672 10968 5681
rect 11020 5672 11022 5681
rect 10966 5607 11022 5616
rect 11072 5234 11100 5782
rect 11256 5710 11284 6072
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11256 5098 11284 5170
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10980 3670 11008 4150
rect 11072 3738 11100 4422
rect 11244 4208 11296 4214
rect 11164 4156 11244 4162
rect 11164 4150 11296 4156
rect 11164 4134 11284 4150
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 11164 3584 11192 4134
rect 11244 3596 11296 3602
rect 11164 3556 11244 3584
rect 10968 3528 11020 3534
rect 10966 3496 10968 3505
rect 11020 3496 11022 3505
rect 11164 3466 11192 3556
rect 11244 3538 11296 3544
rect 10966 3431 11022 3440
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11348 3194 11376 9930
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11440 8974 11468 9658
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11532 7546 11560 11290
rect 11716 11014 11744 11698
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10062 11836 10406
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11624 9654 11652 9930
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11624 8634 11652 9590
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 10612 2746 10824 2774
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10612 2514 10640 2746
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 9048 800 9076 2382
rect 10336 800 10364 2382
rect 11440 1834 11468 7210
rect 11532 5914 11560 7346
rect 11624 6361 11652 8230
rect 11716 8090 11744 9522
rect 11808 8974 11836 9522
rect 11900 9518 11928 11086
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11900 8838 11928 9318
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11716 7954 11744 8026
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11808 7410 11836 7822
rect 11992 7410 12020 11698
rect 12084 8922 12112 13262
rect 12544 12442 12572 17190
rect 12860 17156 13124 17184
rect 12808 17138 12860 17144
rect 12900 17060 12952 17066
rect 12900 17002 12952 17008
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16590 12756 16934
rect 12912 16590 12940 17002
rect 13096 16590 13124 17156
rect 12716 16584 12768 16590
rect 12716 16526 12768 16532
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12912 15570 12940 15914
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 15162 12664 15302
rect 13004 15162 13032 15438
rect 13096 15366 13124 16526
rect 13280 15706 13308 19382
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 13464 16182 13492 16594
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 16182 13584 16390
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13544 16176 13596 16182
rect 13544 16118 13596 16124
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13648 15586 13676 20402
rect 14016 17921 14044 24074
rect 14108 23254 14136 24210
rect 14200 23798 14228 25162
rect 14292 24954 14320 25230
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14292 23610 14320 24890
rect 14568 24614 14596 25842
rect 14832 25832 14884 25838
rect 14832 25774 14884 25780
rect 14844 25702 14872 25774
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14660 24818 14688 25094
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14370 23760 14426 23769
rect 14476 23730 14504 24278
rect 14370 23695 14372 23704
rect 14424 23695 14426 23704
rect 14464 23724 14516 23730
rect 14372 23666 14424 23672
rect 14464 23666 14516 23672
rect 14200 23582 14320 23610
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 14108 23118 14136 23190
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14200 22094 14228 23582
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22166 14320 23054
rect 14384 22710 14412 23122
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14280 22160 14332 22166
rect 14280 22102 14332 22108
rect 14108 22066 14228 22094
rect 14108 19446 14136 22066
rect 14188 22024 14240 22030
rect 14186 21992 14188 22001
rect 14240 21992 14242 22001
rect 14186 21927 14242 21936
rect 14200 21434 14228 21927
rect 14292 21622 14320 22102
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 14476 21865 14504 21966
rect 14462 21856 14518 21865
rect 14462 21791 14518 21800
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14568 21554 14596 24550
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14200 21406 14596 21434
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14200 20369 14228 20402
rect 14186 20360 14242 20369
rect 14384 20330 14412 21014
rect 14186 20295 14242 20304
rect 14372 20324 14424 20330
rect 14372 20266 14424 20272
rect 14476 19530 14504 21286
rect 14568 20602 14596 21406
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14568 19718 14596 20402
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14384 19502 14504 19530
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14200 18834 14228 19314
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14292 18766 14320 19178
rect 14384 18902 14412 19502
rect 14568 19310 14596 19654
rect 14660 19310 14688 24754
rect 14752 24614 14780 24754
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14936 24410 14964 29990
rect 15476 29096 15528 29102
rect 15476 29038 15528 29044
rect 15292 28144 15344 28150
rect 15292 28086 15344 28092
rect 15016 27940 15068 27946
rect 15016 27882 15068 27888
rect 15028 27538 15056 27882
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 15304 27402 15332 28086
rect 15488 27878 15516 29038
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15488 27554 15516 27814
rect 15396 27526 15516 27554
rect 15396 27470 15424 27526
rect 15384 27464 15436 27470
rect 15384 27406 15436 27412
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 15200 26784 15252 26790
rect 15200 26726 15252 26732
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15212 26042 15240 26726
rect 15304 26382 15332 26726
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 15016 25968 15068 25974
rect 15396 25922 15424 27406
rect 15568 27396 15620 27402
rect 15568 27338 15620 27344
rect 15068 25916 15424 25922
rect 15016 25910 15424 25916
rect 15028 25894 15424 25910
rect 15396 24818 15424 25894
rect 15580 24818 15608 27338
rect 15672 25378 15700 29990
rect 15752 29232 15804 29238
rect 15752 29174 15804 29180
rect 15764 28762 15792 29174
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 16120 28144 16172 28150
rect 16120 28086 16172 28092
rect 16132 27674 16160 28086
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16408 27674 16436 27814
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 16396 27668 16448 27674
rect 16396 27610 16448 27616
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15764 26382 15792 26726
rect 15752 26376 15804 26382
rect 15752 26318 15804 26324
rect 15764 26042 15792 26318
rect 15948 26042 15976 26930
rect 16212 26308 16264 26314
rect 16212 26250 16264 26256
rect 16224 26042 16252 26250
rect 16396 26240 16448 26246
rect 16396 26182 16448 26188
rect 15752 26036 15804 26042
rect 15752 25978 15804 25984
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16212 26036 16264 26042
rect 16212 25978 16264 25984
rect 15844 25900 15896 25906
rect 15844 25842 15896 25848
rect 15672 25350 15792 25378
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15568 24812 15620 24818
rect 15568 24754 15620 24760
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 15016 24336 15068 24342
rect 15016 24278 15068 24284
rect 15028 24206 15056 24278
rect 15016 24200 15068 24206
rect 15016 24142 15068 24148
rect 15292 24200 15344 24206
rect 15396 24188 15424 24754
rect 15488 24682 15516 24754
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15568 24200 15620 24206
rect 15344 24160 15516 24188
rect 15292 24142 15344 24148
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14752 22778 14780 22986
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14740 22500 14792 22506
rect 14740 22442 14792 22448
rect 14752 22030 14780 22442
rect 14844 22098 14872 24074
rect 14922 23760 14978 23769
rect 14922 23695 14978 23704
rect 14936 22506 14964 23695
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15120 22982 15148 23598
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 15212 22234 15240 23190
rect 15488 23118 15516 24160
rect 15568 24142 15620 24148
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15396 22506 15424 23054
rect 15488 22778 15516 23054
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15384 22500 15436 22506
rect 15384 22442 15436 22448
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14832 21956 14884 21962
rect 14832 21898 14884 21904
rect 14740 21548 14792 21554
rect 14740 21490 14792 21496
rect 14752 19990 14780 21490
rect 14844 20346 14872 21898
rect 14936 20466 14964 21966
rect 15212 21554 15240 22170
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21690 15332 21830
rect 15292 21684 15344 21690
rect 15292 21626 15344 21632
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15016 20528 15068 20534
rect 15016 20470 15068 20476
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14844 20318 14964 20346
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14936 19854 14964 20318
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 15028 19786 15056 20470
rect 15108 20460 15160 20466
rect 15396 20448 15424 21966
rect 15580 21690 15608 24142
rect 15672 22030 15700 24142
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15488 21078 15516 21490
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15580 21146 15608 21422
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15476 21072 15528 21078
rect 15476 21014 15528 21020
rect 15160 20420 15424 20448
rect 15108 20402 15160 20408
rect 15120 19854 15148 20402
rect 15488 19938 15516 21014
rect 15488 19910 15608 19938
rect 15580 19854 15608 19910
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 15028 19378 15056 19722
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 14556 19304 14608 19310
rect 14648 19304 14700 19310
rect 14556 19246 14608 19252
rect 14646 19272 14648 19281
rect 14700 19272 14702 19281
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14384 18766 14412 18838
rect 14568 18766 14596 19246
rect 14646 19207 14702 19216
rect 14752 18766 14780 19314
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14002 17912 14058 17921
rect 14002 17847 14058 17856
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13740 17202 13768 17750
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13740 16522 13768 17138
rect 14292 17134 14320 18226
rect 14936 18154 14964 18566
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 15120 17542 15148 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15212 18358 15240 19450
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 18698 15332 19110
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15304 18426 15332 18634
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15200 18352 15252 18358
rect 15200 18294 15252 18300
rect 15660 18080 15712 18086
rect 15660 18022 15712 18028
rect 15672 17678 15700 18022
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13740 16250 13768 16458
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13556 15558 13676 15586
rect 14016 15570 14044 17070
rect 14292 16590 14320 17070
rect 14648 16720 14700 16726
rect 14648 16662 14700 16668
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16182 14320 16390
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14004 15564 14056 15570
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14414 13124 14894
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12992 14340 13044 14346
rect 12992 14282 13044 14288
rect 13004 13938 13032 14282
rect 13096 14006 13124 14350
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 11801 12664 13670
rect 12820 13326 12848 13670
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12912 12238 12940 13126
rect 13096 12714 13124 13806
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 12622 11792 12678 11801
rect 12912 11762 12940 12174
rect 13004 11762 13032 12174
rect 12622 11727 12678 11736
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 12716 11688 12768 11694
rect 12714 11656 12716 11665
rect 12808 11688 12860 11694
rect 12768 11656 12770 11665
rect 12808 11630 12860 11636
rect 12714 11591 12770 11600
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 12268 10470 12296 11154
rect 12544 11150 12572 11494
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10742 12480 11018
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12440 10736 12492 10742
rect 12440 10678 12492 10684
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 9042 12204 9318
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12084 8894 12204 8922
rect 12176 7818 12204 8894
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12440 8492 12492 8498
rect 12440 8434 12492 8440
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11716 6662 11744 7346
rect 11808 6730 11836 7346
rect 12084 6798 12112 7754
rect 12360 7410 12388 8434
rect 12452 8294 12480 8434
rect 12544 8430 12572 10950
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12636 8090 12664 9998
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12636 7478 12664 8026
rect 12728 7546 12756 11086
rect 12820 10266 12848 11630
rect 13096 11626 13124 12174
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12912 11393 12940 11494
rect 12898 11384 12954 11393
rect 12898 11319 12954 11328
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12912 10810 12940 11154
rect 13004 11014 13032 11494
rect 13082 11384 13138 11393
rect 13082 11319 13138 11328
rect 13096 11014 13124 11319
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13084 11008 13136 11014
rect 13084 10950 13136 10956
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12912 10198 12940 10746
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13096 9994 13124 10610
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13096 9518 13124 9930
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13004 8974 13032 9386
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12820 8634 12848 8910
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12912 7546 12940 8910
rect 13096 8616 13124 9454
rect 13188 9178 13216 15438
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14822 13308 14962
rect 13556 14890 13584 15558
rect 14004 15506 14056 15512
rect 14292 15366 14320 15982
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13372 13938 13400 14758
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13268 12368 13320 12374
rect 13268 12310 13320 12316
rect 13280 11642 13308 12310
rect 13372 11778 13400 13874
rect 13464 13326 13492 14214
rect 13648 13938 13676 14214
rect 13832 14006 13860 14350
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 14016 13938 14044 14418
rect 14108 13938 14136 14826
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14200 14482 14228 14554
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13544 13864 13596 13870
rect 14108 13841 14136 13874
rect 13544 13806 13596 13812
rect 14094 13832 14150 13841
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13556 12238 13584 13806
rect 14094 13767 14150 13776
rect 14292 13394 14320 14894
rect 14384 14414 14412 15438
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 14618 14596 14894
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14660 14414 14688 16662
rect 15028 14482 15056 17070
rect 15304 15570 15332 17478
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15488 16250 15516 16458
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15570 15700 15846
rect 15292 15564 15344 15570
rect 15212 15524 15292 15552
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14568 14006 14596 14282
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14660 13802 14688 14350
rect 15028 14346 15056 14418
rect 15212 14414 15240 15524
rect 15292 15506 15344 15512
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12850 14320 13330
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13372 11762 13584 11778
rect 13372 11756 13596 11762
rect 13372 11750 13544 11756
rect 13544 11698 13596 11704
rect 13280 11614 13400 11642
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13280 10742 13308 11154
rect 13372 10742 13400 11614
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 10062 13308 10134
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13280 9654 13308 9998
rect 13268 9648 13320 9654
rect 13268 9590 13320 9596
rect 13556 9586 13584 11698
rect 13648 11694 13676 12650
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 14188 12164 14240 12170
rect 13832 12102 13860 12135
rect 14188 12106 14240 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 13636 11688 13688 11694
rect 13924 11665 13952 11698
rect 13636 11630 13688 11636
rect 13910 11656 13966 11665
rect 13728 11620 13780 11626
rect 13910 11591 13966 11600
rect 13728 11562 13780 11568
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13648 10198 13676 10610
rect 13740 10266 13768 11562
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13924 10742 13952 11086
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13740 9722 13768 10202
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 13096 8588 13308 8616
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12360 6866 12388 7346
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12360 6730 12388 6802
rect 12452 6798 12480 7278
rect 12820 7002 12848 7278
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11610 6352 11666 6361
rect 11716 6322 11744 6598
rect 11808 6390 11836 6666
rect 12636 6458 12664 6734
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11610 6287 11666 6296
rect 11704 6316 11756 6322
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11624 5778 11652 6287
rect 11704 6258 11756 6264
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11716 5710 11744 6054
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11808 5250 11836 6054
rect 11624 5234 11836 5250
rect 11612 5228 11836 5234
rect 11664 5222 11836 5228
rect 11612 5170 11664 5176
rect 11900 5030 11928 6326
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5370 12020 5646
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12084 5234 12112 6258
rect 12636 5710 12664 6394
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 11612 4480 11664 4486
rect 11532 4440 11612 4468
rect 11532 2922 11560 4440
rect 11612 4422 11664 4428
rect 11716 4128 11744 4558
rect 11900 4282 11928 4558
rect 11992 4554 12020 5170
rect 12084 4758 12112 5170
rect 12072 4752 12124 4758
rect 12072 4694 12124 4700
rect 12728 4622 12756 6802
rect 12912 6458 12940 7346
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13004 5692 13032 8434
rect 13280 7868 13308 8588
rect 13740 8430 13768 9522
rect 13832 8650 13860 10406
rect 14016 9994 14044 12038
rect 14200 11762 14228 12106
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14094 11656 14150 11665
rect 14094 11591 14150 11600
rect 14108 10810 14136 11591
rect 14292 11150 14320 12786
rect 14844 12442 14872 12854
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14936 12238 14964 12582
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11830 14596 12038
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14844 11665 14872 11698
rect 14830 11656 14886 11665
rect 14830 11591 14886 11600
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 11354 14780 11494
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14292 10130 14320 11086
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13832 8634 13952 8650
rect 13820 8628 13952 8634
rect 13872 8622 13952 8628
rect 13820 8570 13872 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13464 7886 13492 8366
rect 13832 8090 13860 8434
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13726 7984 13782 7993
rect 13832 7954 13860 8026
rect 13726 7919 13782 7928
rect 13820 7948 13872 7954
rect 13740 7886 13768 7919
rect 13820 7890 13872 7896
rect 13924 7886 13952 8622
rect 14292 8498 14320 10066
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13452 7880 13504 7886
rect 13280 7840 13400 7868
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13096 6866 13124 7482
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13280 6798 13308 7239
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13084 5704 13136 5710
rect 13004 5672 13084 5692
rect 13136 5672 13138 5681
rect 13004 5664 13082 5672
rect 13280 5642 13308 6734
rect 13082 5607 13138 5616
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13084 5228 13136 5234
rect 13188 5216 13216 5578
rect 13268 5228 13320 5234
rect 13188 5188 13268 5216
rect 13084 5170 13136 5176
rect 13268 5170 13320 5176
rect 13096 5098 13124 5170
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13096 4826 13124 5034
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13280 4622 13308 5170
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 12268 4214 12296 4490
rect 12636 4214 12664 4558
rect 12728 4282 12756 4558
rect 13280 4282 13308 4558
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 11796 4140 11848 4146
rect 11716 4100 11796 4128
rect 11796 4082 11848 4088
rect 12728 3738 12756 4218
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13188 4010 13216 4082
rect 13176 4004 13228 4010
rect 13096 3964 13176 3992
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 13096 3534 13124 3964
rect 13176 3946 13228 3952
rect 13372 3942 13400 7840
rect 13452 7822 13504 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13556 7410 13584 7686
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 6322 13768 7278
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13464 5166 13492 5646
rect 13542 5264 13598 5273
rect 13542 5199 13544 5208
rect 13596 5199 13598 5208
rect 13740 5216 13768 6258
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13832 5914 13860 6190
rect 13924 5914 13952 6258
rect 14016 5953 14044 7346
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6322 14136 6598
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14002 5944 14058 5953
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13912 5908 13964 5914
rect 14002 5879 14058 5888
rect 13912 5850 13964 5856
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13832 5370 13860 5646
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13820 5228 13872 5234
rect 13740 5188 13820 5216
rect 13544 5170 13596 5176
rect 13820 5170 13872 5176
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13556 4690 13584 5170
rect 14016 5166 14044 5879
rect 14096 5364 14148 5370
rect 14200 5352 14228 7822
rect 14148 5324 14228 5352
rect 14096 5306 14148 5312
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13084 3528 13136 3534
rect 12162 3496 12218 3505
rect 11980 3460 12032 3466
rect 13084 3470 13136 3476
rect 12162 3431 12218 3440
rect 11980 3402 12032 3408
rect 11992 3194 12020 3402
rect 12176 3194 12204 3431
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 13280 3126 13308 3674
rect 13464 3534 13492 4082
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 3738 13676 4014
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13832 3466 13860 4150
rect 13820 3460 13872 3466
rect 13820 3402 13872 3408
rect 11704 3120 11756 3126
rect 13268 3120 13320 3126
rect 11756 3080 11928 3108
rect 11704 3062 11756 3068
rect 11900 3074 11928 3080
rect 11900 3058 12112 3074
rect 13268 3062 13320 3068
rect 11900 3052 12124 3058
rect 11900 3046 12072 3052
rect 12072 2994 12124 3000
rect 11612 2984 11664 2990
rect 11664 2944 12020 2972
rect 11612 2926 11664 2932
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 11992 2854 12020 2944
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11900 2514 11928 2790
rect 12070 2680 12126 2689
rect 12070 2615 12072 2624
rect 12124 2615 12126 2624
rect 12808 2644 12860 2650
rect 12072 2586 12124 2592
rect 12808 2586 12860 2592
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 12820 2446 12848 2586
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 11428 1828 11480 1834
rect 11428 1770 11480 1776
rect 11624 800 11652 2314
rect 12912 800 12940 2382
rect 13280 1902 13308 2382
rect 14016 2038 14044 5102
rect 14292 3602 14320 8434
rect 14384 7970 14412 9930
rect 14384 7942 14596 7970
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14384 7546 14412 7822
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14476 7410 14504 7822
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 4826 14412 5170
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3194 14320 3538
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14004 2032 14056 2038
rect 14004 1974 14056 1980
rect 13268 1896 13320 1902
rect 13268 1838 13320 1844
rect 14200 800 14228 2314
rect 14476 1698 14504 7346
rect 14568 4214 14596 7942
rect 14660 7886 14688 10746
rect 14936 10742 14964 12174
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 15028 11626 15056 11727
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 15028 10674 15056 11290
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14936 9654 14964 9930
rect 14924 9648 14976 9654
rect 15304 9625 15332 15370
rect 15672 14414 15700 15506
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 13394 15700 13670
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15764 12306 15792 25350
rect 15856 25294 15884 25842
rect 16224 25838 16252 25978
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16408 25702 16436 26182
rect 16396 25696 16448 25702
rect 16396 25638 16448 25644
rect 15844 25288 15896 25294
rect 15844 25230 15896 25236
rect 15856 24954 15884 25230
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 15948 24886 15976 25094
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 16592 24614 16620 30126
rect 20720 30116 20772 30122
rect 20720 30058 20772 30064
rect 22376 30116 22428 30122
rect 22376 30058 22428 30064
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 19524 30048 19576 30054
rect 19524 29990 19576 29996
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 17880 28558 17908 29242
rect 18052 29096 18104 29102
rect 18052 29038 18104 29044
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 17408 28552 17460 28558
rect 17408 28494 17460 28500
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16776 27402 16804 27814
rect 16960 27470 16988 28494
rect 17420 28218 17448 28494
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17604 28218 17632 28358
rect 17408 28212 17460 28218
rect 17408 28154 17460 28160
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17144 27606 17172 28018
rect 17604 27606 17632 28154
rect 17868 27872 17920 27878
rect 17868 27814 17920 27820
rect 17880 27674 17908 27814
rect 17868 27668 17920 27674
rect 17868 27610 17920 27616
rect 17132 27600 17184 27606
rect 17132 27542 17184 27548
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16868 26586 17172 26602
rect 16856 26580 17172 26586
rect 16908 26574 17172 26580
rect 16856 26522 16908 26528
rect 17144 26518 17172 26574
rect 17132 26512 17184 26518
rect 16868 26438 17080 26466
rect 17132 26454 17184 26460
rect 16868 25906 16896 26438
rect 17052 26382 17080 26438
rect 17224 26444 17276 26450
rect 17224 26386 17276 26392
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16684 24954 16712 25230
rect 16868 24954 16896 25842
rect 16960 25498 16988 26318
rect 17236 26296 17264 26386
rect 17684 26308 17736 26314
rect 17236 26268 17684 26296
rect 17788 26296 17816 27542
rect 17972 27402 18000 28358
rect 18064 27674 18092 29038
rect 18236 28552 18288 28558
rect 18236 28494 18288 28500
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17868 26852 17920 26858
rect 17868 26794 17920 26800
rect 17736 26268 17816 26296
rect 17684 26250 17736 26256
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 17684 25968 17736 25974
rect 17684 25910 17736 25916
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 17052 25430 17080 25910
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17040 25424 17092 25430
rect 17040 25366 17092 25372
rect 17040 25288 17092 25294
rect 17144 25276 17172 25842
rect 17592 25832 17644 25838
rect 17592 25774 17644 25780
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17420 25294 17448 25638
rect 17604 25498 17632 25774
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 17092 25248 17172 25276
rect 17408 25288 17460 25294
rect 17406 25256 17408 25265
rect 17460 25256 17462 25265
rect 17040 25230 17092 25236
rect 16672 24948 16724 24954
rect 16672 24890 16724 24896
rect 16856 24948 16908 24954
rect 16856 24890 16908 24896
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16960 24682 16988 24754
rect 16948 24676 17000 24682
rect 16948 24618 17000 24624
rect 16580 24608 16632 24614
rect 17052 24585 17080 25230
rect 17406 25191 17462 25200
rect 17328 24818 17448 24834
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17316 24812 17448 24818
rect 17368 24806 17448 24812
rect 17316 24754 17368 24760
rect 16580 24550 16632 24556
rect 17038 24576 17094 24585
rect 17038 24511 17094 24520
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 16868 24206 16896 24346
rect 16960 24206 16988 24346
rect 15844 24200 15896 24206
rect 16856 24200 16908 24206
rect 15844 24142 15896 24148
rect 16776 24160 16856 24188
rect 15856 23798 15884 24142
rect 16672 24064 16724 24070
rect 16672 24006 16724 24012
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 16684 23322 16712 24006
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16408 22778 16436 23054
rect 16684 22982 16712 23054
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16396 22772 16448 22778
rect 16396 22714 16448 22720
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16132 20369 16160 22578
rect 16776 22030 16804 24160
rect 16856 24142 16908 24148
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 17040 24132 17092 24138
rect 17040 24074 17092 24080
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23526 16988 24006
rect 17052 23730 17080 24074
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16868 23050 16896 23462
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16960 23050 16988 23258
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 16868 22710 16896 22986
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16960 22545 16988 22578
rect 16946 22536 17002 22545
rect 16946 22471 17002 22480
rect 17144 22094 17172 24754
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17236 23798 17264 24142
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 17328 23610 17356 24618
rect 17420 24410 17448 24806
rect 17500 24812 17552 24818
rect 17500 24754 17552 24760
rect 17512 24682 17540 24754
rect 17696 24698 17724 25910
rect 17788 24818 17816 26268
rect 17880 25906 17908 26794
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18064 25906 18092 26318
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 18156 25906 18184 26250
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 17868 25356 17920 25362
rect 17868 25298 17920 25304
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17500 24676 17552 24682
rect 17696 24670 17816 24698
rect 17500 24618 17552 24624
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 16960 22066 17172 22094
rect 17236 23582 17356 23610
rect 16764 22024 16816 22030
rect 16764 21966 16816 21972
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16304 21344 16356 21350
rect 16304 21286 16356 21292
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 20466 16252 20810
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16316 20380 16344 21286
rect 16408 20942 16436 21558
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16868 21457 16896 21490
rect 16854 21448 16910 21457
rect 16854 21383 16910 21392
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16396 20392 16448 20398
rect 16118 20360 16174 20369
rect 16316 20352 16396 20380
rect 16396 20334 16448 20340
rect 16118 20295 16174 20304
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16224 19990 16252 20198
rect 16212 19984 16264 19990
rect 16212 19926 16264 19932
rect 16028 19236 16080 19242
rect 16028 19178 16080 19184
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18766 15884 19110
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15856 18290 15884 18702
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15948 14618 15976 16050
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16040 13938 16068 19178
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 14498 16160 15982
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16316 15094 16344 15438
rect 16212 15088 16264 15094
rect 16212 15030 16264 15036
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16224 14618 16252 15030
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16132 14470 16252 14498
rect 16408 14482 16436 15846
rect 16500 15706 16528 20946
rect 16592 20942 16620 21286
rect 16580 20936 16632 20942
rect 16960 20890 16988 22066
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17040 21412 17092 21418
rect 17040 21354 17092 21360
rect 17052 20942 17080 21354
rect 17144 21350 17172 21966
rect 17236 21894 17264 23582
rect 17420 22778 17448 24142
rect 17512 23848 17540 24618
rect 17592 24608 17644 24614
rect 17684 24608 17736 24614
rect 17592 24550 17644 24556
rect 17682 24576 17684 24585
rect 17736 24576 17738 24585
rect 17604 24410 17632 24550
rect 17682 24511 17738 24520
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 17604 24206 17632 24346
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17512 23820 17632 23848
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17316 22704 17368 22710
rect 17316 22646 17368 22652
rect 17328 22234 17356 22646
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17328 21554 17356 22170
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17236 21010 17264 21490
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 16580 20878 16632 20884
rect 16776 20862 16988 20890
rect 17040 20936 17092 20942
rect 17040 20878 17092 20884
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 20466 16712 20742
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16776 20058 16804 20862
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16868 20466 16896 20742
rect 16856 20460 16908 20466
rect 16856 20402 16908 20408
rect 16960 20262 16988 20742
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17040 20392 17092 20398
rect 17038 20360 17040 20369
rect 17092 20360 17094 20369
rect 17038 20295 17094 20304
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16684 19786 16712 19994
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16590 16620 16934
rect 16684 16658 16712 19722
rect 16776 19310 16804 19994
rect 16960 19378 16988 19994
rect 17052 19553 17080 20295
rect 17144 19990 17172 20402
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17038 19544 17094 19553
rect 17144 19514 17172 19926
rect 17038 19479 17094 19488
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16868 18970 16896 19314
rect 16960 19242 16988 19314
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 17144 18902 17172 19450
rect 17132 18896 17184 18902
rect 17132 18838 17184 18844
rect 17236 18850 17264 20946
rect 17328 20058 17356 21286
rect 17316 20052 17368 20058
rect 17316 19994 17368 20000
rect 17420 19938 17448 21830
rect 17512 21457 17540 23666
rect 17498 21448 17554 21457
rect 17498 21383 17554 21392
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17328 19910 17448 19938
rect 17328 19446 17356 19910
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17144 18766 17172 18838
rect 17236 18822 17356 18850
rect 17328 18766 17356 18822
rect 17420 18766 17448 19790
rect 17512 19786 17540 20266
rect 17604 19854 17632 23820
rect 17696 22642 17724 24511
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17684 21548 17736 21554
rect 17684 21490 17736 21496
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17696 19394 17724 21490
rect 17512 19378 17724 19394
rect 17500 19372 17724 19378
rect 17552 19366 17724 19372
rect 17500 19314 17552 19320
rect 17682 18864 17738 18873
rect 17788 18834 17816 24670
rect 17880 22692 17908 25298
rect 17960 24880 18012 24886
rect 18012 24840 18092 24868
rect 17960 24822 18012 24828
rect 18064 24585 18092 24840
rect 18050 24576 18106 24585
rect 18050 24511 18106 24520
rect 18064 24206 18092 24511
rect 18248 24410 18276 28494
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 17972 23118 18000 23802
rect 18156 23798 18184 24006
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 18340 23322 18368 29990
rect 18788 29232 18840 29238
rect 18788 29174 18840 29180
rect 18512 28960 18564 28966
rect 18512 28902 18564 28908
rect 18524 28626 18552 28902
rect 18800 28762 18828 29174
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18512 28620 18564 28626
rect 18512 28562 18564 28568
rect 18524 28082 18552 28562
rect 19248 28212 19300 28218
rect 19248 28154 19300 28160
rect 18512 28076 18564 28082
rect 18512 28018 18564 28024
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 27674 19012 28018
rect 18972 27668 19024 27674
rect 18972 27610 19024 27616
rect 19260 27470 19288 28154
rect 19432 28144 19484 28150
rect 19432 28086 19484 28092
rect 19444 27878 19472 28086
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19444 27674 19472 27814
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19352 27130 19380 27270
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 18420 26852 18472 26858
rect 18420 26794 18472 26800
rect 18432 26382 18460 26794
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18432 25498 18460 25842
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18524 25378 18552 27066
rect 19248 27056 19300 27062
rect 19248 26998 19300 27004
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18616 26382 18644 26930
rect 18708 26382 18736 26930
rect 19260 26382 19288 26998
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18972 26376 19024 26382
rect 18972 26318 19024 26324
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 18616 26042 18644 26318
rect 18788 26308 18840 26314
rect 18788 26250 18840 26256
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18800 25770 18828 26250
rect 18984 25974 19012 26318
rect 19352 26246 19380 27066
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 19444 25974 19472 27610
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 18788 25764 18840 25770
rect 18788 25706 18840 25712
rect 19432 25764 19484 25770
rect 19432 25706 19484 25712
rect 18524 25350 18644 25378
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18420 24812 18472 24818
rect 18420 24754 18472 24760
rect 18432 24342 18460 24754
rect 18420 24336 18472 24342
rect 18420 24278 18472 24284
rect 18432 24206 18460 24278
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18328 23316 18380 23322
rect 18248 23276 18328 23304
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 18064 22778 18092 23054
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22704 18012 22710
rect 17880 22664 17960 22692
rect 17960 22646 18012 22652
rect 17868 22568 17920 22574
rect 17866 22536 17868 22545
rect 17920 22536 17922 22545
rect 17866 22471 17922 22480
rect 18248 21026 18276 23276
rect 18328 23258 18380 23264
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18340 22710 18368 23054
rect 18328 22704 18380 22710
rect 18328 22646 18380 22652
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18248 20998 18368 21026
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19854 17908 20198
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17972 19786 18000 20878
rect 18064 20466 18092 20878
rect 18236 20868 18288 20874
rect 18236 20810 18288 20816
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 18064 19990 18092 20402
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18156 20058 18184 20334
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18052 19984 18104 19990
rect 18248 19938 18276 20810
rect 18340 20466 18368 20998
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18052 19926 18104 19932
rect 18156 19910 18276 19938
rect 18156 19854 18184 19910
rect 18340 19854 18368 20402
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17866 19544 17922 19553
rect 17866 19479 17922 19488
rect 17880 19446 17908 19479
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17960 19440 18012 19446
rect 17960 19382 18012 19388
rect 17682 18799 17738 18808
rect 17776 18828 17828 18834
rect 17696 18766 17724 18799
rect 17776 18770 17828 18776
rect 17972 18766 18000 19382
rect 18156 18970 18184 19790
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18248 19514 18276 19722
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18328 19372 18380 19378
rect 18432 19360 18460 22578
rect 18380 19332 18460 19360
rect 18328 19314 18380 19320
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16776 18290 16804 18566
rect 16868 18358 16896 18566
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 17052 18290 17080 18566
rect 17512 18426 17540 18702
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17696 18290 17724 18702
rect 17972 18290 18000 18702
rect 18340 18698 18368 19314
rect 18328 18692 18380 18698
rect 18328 18634 18380 18640
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18340 18290 18368 18362
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 17696 18154 17724 18226
rect 16856 18148 16908 18154
rect 16856 18090 16908 18096
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16040 13394 16068 13874
rect 16224 13870 16252 14470
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15856 12442 15884 12854
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 16224 12306 16252 13806
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 14924 9590 14976 9596
rect 15290 9616 15346 9625
rect 15290 9551 15346 9560
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15580 8974 15608 9318
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15568 8968 15620 8974
rect 15568 8910 15620 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8566 14780 8774
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15488 8090 15516 8502
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7478 14688 7822
rect 15672 7546 15700 8978
rect 16224 8838 16252 9998
rect 16408 9042 16436 12242
rect 16500 11830 16528 15642
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13258 16804 13670
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16488 11824 16540 11830
rect 16488 11766 16540 11772
rect 16500 11218 16528 11766
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16684 11150 16712 12174
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16684 9586 16712 11086
rect 16762 10704 16818 10713
rect 16762 10639 16764 10648
rect 16816 10639 16818 10648
rect 16764 10610 16816 10616
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8634 16252 8774
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15304 7002 15332 7278
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15028 6361 15056 6802
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15014 6352 15070 6361
rect 14648 6316 14700 6322
rect 14700 6276 14780 6304
rect 15014 6287 15016 6296
rect 14648 6258 14700 6264
rect 14648 5704 14700 5710
rect 14648 5646 14700 5652
rect 14660 5370 14688 5646
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14752 4622 14780 6276
rect 15068 6287 15070 6296
rect 15016 6258 15068 6264
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4826 14872 5170
rect 14936 4826 14964 6054
rect 15212 5250 15240 6598
rect 15120 5234 15240 5250
rect 15108 5228 15240 5234
rect 15160 5222 15240 5228
rect 15108 5170 15160 5176
rect 15016 5160 15068 5166
rect 15016 5102 15068 5108
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14740 4616 14792 4622
rect 15028 4604 15056 5102
rect 15108 4616 15160 4622
rect 15028 4576 15108 4604
rect 14740 4558 14792 4564
rect 15108 4558 15160 4564
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14660 3602 14688 3946
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14752 3194 14780 3878
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14844 3074 14872 4082
rect 15304 3602 15332 6666
rect 15580 6254 15608 6734
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 6322 15700 6598
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15384 6248 15436 6254
rect 15384 6190 15436 6196
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15396 5098 15424 6190
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15488 5234 15516 5782
rect 15764 5710 15792 6802
rect 16132 6798 16160 8502
rect 16408 8430 16436 8978
rect 16684 8838 16712 9522
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16684 7886 16712 8774
rect 16776 8401 16804 10610
rect 16762 8392 16818 8401
rect 16762 8327 16818 8336
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 15752 5704 15804 5710
rect 15750 5672 15752 5681
rect 15804 5672 15806 5681
rect 15660 5636 15712 5642
rect 15750 5607 15806 5616
rect 15660 5578 15712 5584
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15488 4622 15516 5170
rect 15580 4826 15608 5170
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15488 4282 15516 4558
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15396 3194 15424 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 14752 3046 14872 3074
rect 14752 2854 14780 3046
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 14464 1692 14516 1698
rect 14464 1634 14516 1640
rect 15488 800 15516 2314
rect 15580 2310 15608 4762
rect 15672 2310 15700 5578
rect 16224 5234 16252 6734
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16500 5370 16528 5850
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16132 5098 16160 5170
rect 16120 5092 16172 5098
rect 16120 5034 16172 5040
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16132 3126 16160 3334
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16224 2650 16252 5170
rect 16592 4826 16620 7346
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16684 5914 16712 6666
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16776 5234 16804 6802
rect 16868 5794 16896 18090
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17328 17746 17356 18022
rect 18340 17882 18368 18226
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17316 17740 17368 17746
rect 17316 17682 17368 17688
rect 17972 16794 18000 17750
rect 18432 17678 18460 18226
rect 18524 18086 18552 25230
rect 18616 18426 18644 25350
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18892 23526 18920 24754
rect 18984 24585 19012 24754
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 18970 24576 19026 24585
rect 18970 24511 19026 24520
rect 19168 23662 19196 24618
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19352 24274 19380 24346
rect 19340 24268 19392 24274
rect 19340 24210 19392 24216
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19260 23866 19288 24074
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 19156 23316 19208 23322
rect 19156 23258 19208 23264
rect 19064 23248 19116 23254
rect 19064 23190 19116 23196
rect 18696 23112 18748 23118
rect 18696 23054 18748 23060
rect 18708 22506 18736 23054
rect 18696 22500 18748 22506
rect 18696 22442 18748 22448
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18800 21078 18828 21490
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18892 20754 18920 22442
rect 19076 22438 19104 23190
rect 19168 22642 19196 23258
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 19352 22030 19380 24210
rect 19444 23118 19472 25706
rect 19536 25158 19564 29990
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 19616 27600 19668 27606
rect 19616 27542 19668 27548
rect 19628 26382 19656 27542
rect 19996 27538 20024 28562
rect 20260 28484 20312 28490
rect 20260 28426 20312 28432
rect 20272 28218 20300 28426
rect 20260 28212 20312 28218
rect 20260 28154 20312 28160
rect 19984 27532 20036 27538
rect 19984 27474 20036 27480
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19720 25362 19748 27406
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19812 25906 19840 26182
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19892 25900 19944 25906
rect 19996 25888 20024 27474
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 27130 20668 27270
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 19944 25860 20024 25888
rect 19892 25842 19944 25848
rect 19708 25356 19760 25362
rect 19708 25298 19760 25304
rect 19524 25152 19576 25158
rect 19524 25094 19576 25100
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19536 23866 19564 24754
rect 19720 24682 19748 25298
rect 19800 25152 19852 25158
rect 19800 25094 19852 25100
rect 19708 24676 19760 24682
rect 19708 24618 19760 24624
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19706 24576 19762 24585
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19444 22710 19472 23054
rect 19432 22704 19484 22710
rect 19432 22646 19484 22652
rect 19536 22098 19564 23802
rect 19628 23730 19656 24550
rect 19706 24511 19762 24520
rect 19720 24206 19748 24511
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19708 24064 19760 24070
rect 19708 24006 19760 24012
rect 19720 23866 19748 24006
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19812 23610 19840 25094
rect 19996 24818 20024 25860
rect 20088 25294 20116 26318
rect 20260 26308 20312 26314
rect 20260 26250 20312 26256
rect 20272 25974 20300 26250
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20536 25356 20588 25362
rect 20536 25298 20588 25304
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 20088 24682 20116 24822
rect 20076 24676 20128 24682
rect 20076 24618 20128 24624
rect 19984 24336 20036 24342
rect 19984 24278 20036 24284
rect 19996 24120 20024 24278
rect 20548 24256 20576 25298
rect 20640 24682 20668 27066
rect 20732 26858 20760 30058
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 21100 28422 21128 29106
rect 21272 28484 21324 28490
rect 21272 28426 21324 28432
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 21100 28014 21128 28358
rect 21284 28218 21312 28426
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 22020 28150 22048 28426
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 21088 28008 21140 28014
rect 21088 27950 21140 27956
rect 21100 26994 21128 27950
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21192 27130 21220 27338
rect 21180 27124 21232 27130
rect 21180 27066 21232 27072
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 21824 26240 21876 26246
rect 21824 26182 21876 26188
rect 21836 26042 21864 26182
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21468 25498 21496 25910
rect 22020 25838 22048 26930
rect 22284 25968 22336 25974
rect 22284 25910 22336 25916
rect 22008 25832 22060 25838
rect 22008 25774 22060 25780
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 22020 25294 22048 25774
rect 22296 25498 22324 25910
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 21272 24948 21324 24954
rect 21272 24890 21324 24896
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20548 24228 20668 24256
rect 20536 24194 20588 24200
rect 20076 24132 20128 24138
rect 20536 24136 20588 24142
rect 19996 24092 20076 24120
rect 20076 24074 20128 24080
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23798 19932 24006
rect 19892 23792 19944 23798
rect 19892 23734 19944 23740
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19720 23582 19840 23610
rect 19720 22778 19748 23582
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19892 23520 19944 23526
rect 19892 23462 19944 23468
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19720 22642 19748 22714
rect 19812 22642 19840 23462
rect 19708 22636 19760 22642
rect 19708 22578 19760 22584
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19340 22024 19392 22030
rect 19154 21992 19210 22001
rect 19340 21966 19392 21972
rect 19154 21927 19156 21936
rect 19208 21927 19210 21936
rect 19156 21898 19208 21904
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19076 21350 19104 21490
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 21010 19104 21286
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 18800 20726 18920 20754
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18708 19854 18736 20402
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18800 19786 18828 20726
rect 19352 20466 19380 21830
rect 19536 21554 19564 22034
rect 19720 22030 19748 22578
rect 19904 22574 19932 23462
rect 19996 22642 20024 23666
rect 20548 23526 20576 24136
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20168 22704 20220 22710
rect 20168 22646 20220 22652
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19996 22234 20024 22578
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19892 21956 19944 21962
rect 19892 21898 19944 21904
rect 19524 21548 19576 21554
rect 19524 21490 19576 21496
rect 19536 20942 19564 21490
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19444 20602 19472 20878
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19524 20460 19576 20466
rect 19628 20448 19656 21286
rect 19576 20420 19748 20448
rect 19524 20402 19576 20408
rect 19340 20324 19392 20330
rect 19524 20324 19576 20330
rect 19392 20284 19524 20312
rect 19340 20266 19392 20272
rect 19524 20266 19576 20272
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18800 19360 18828 19722
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18708 19332 18828 19360
rect 18708 18970 18736 19332
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18708 17814 18736 18906
rect 18892 18902 18920 19382
rect 18984 19378 19012 19790
rect 19260 19786 19288 19887
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19260 19360 19288 19722
rect 19444 19446 19472 19994
rect 19616 19848 19668 19854
rect 19522 19816 19578 19825
rect 19616 19790 19668 19796
rect 19522 19751 19578 19760
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19340 19372 19392 19378
rect 19260 19332 19340 19360
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18984 18766 19012 19314
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 18170 18920 18634
rect 18984 18290 19012 18702
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18892 18142 19012 18170
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18432 17270 18460 17614
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16794 18184 17070
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 17408 16720 17460 16726
rect 17408 16662 17460 16668
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17420 16590 17448 16662
rect 18064 16590 18092 16662
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 15162 17356 15438
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17420 15026 17448 16526
rect 17880 16454 17908 16526
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17512 15978 17540 16390
rect 17788 16182 17816 16390
rect 17776 16176 17828 16182
rect 17776 16118 17828 16124
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17512 15502 17540 15914
rect 17604 15502 17632 15982
rect 17788 15570 17816 16118
rect 17880 16046 17908 16390
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17972 15978 18000 16526
rect 18064 16028 18092 16526
rect 18144 16040 18196 16046
rect 18064 16000 18144 16028
rect 18144 15982 18196 15988
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 18248 15706 18276 17138
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17972 14550 18000 15506
rect 18236 15428 18288 15434
rect 18236 15370 18288 15376
rect 18248 14822 18276 15370
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18248 14550 18276 14758
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 18236 14544 18288 14550
rect 18512 14544 18564 14550
rect 18236 14486 18288 14492
rect 18326 14512 18382 14521
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17052 13938 17080 14282
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17052 13308 17080 13874
rect 17420 13870 17448 14214
rect 18156 13938 18184 14350
rect 18248 14278 18276 14486
rect 18512 14486 18564 14492
rect 18602 14512 18658 14521
rect 18326 14447 18328 14456
rect 18380 14447 18382 14456
rect 18328 14418 18380 14424
rect 18524 14414 18552 14486
rect 18602 14447 18604 14456
rect 18656 14447 18658 14456
rect 18604 14418 18656 14424
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18340 14074 18368 14282
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18708 13938 18736 16186
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 18236 13932 18288 13938
rect 18236 13874 18288 13880
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 18248 13394 18276 13874
rect 18708 13394 18736 13874
rect 18236 13388 18288 13394
rect 18236 13330 18288 13336
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 17132 13320 17184 13326
rect 17052 13280 17132 13308
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16960 12442 16988 12718
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17052 12238 17080 13280
rect 17132 13262 17184 13268
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17696 12918 17724 13126
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17880 12102 17908 12922
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17512 11898 17540 12038
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17236 11286 17264 11630
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 17052 10606 17080 11086
rect 17328 11014 17356 11698
rect 17880 11150 17908 12038
rect 17592 11144 17644 11150
rect 17512 11104 17592 11132
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17052 9586 17080 10202
rect 17328 9994 17356 10950
rect 17420 10674 17448 10950
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17408 10464 17460 10470
rect 17408 10406 17460 10412
rect 17316 9988 17368 9994
rect 17316 9930 17368 9936
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16960 9178 16988 9454
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 17420 8974 17448 10406
rect 17512 10130 17540 11104
rect 17592 11086 17644 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17880 10674 17908 11086
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 10198 17908 10610
rect 17868 10192 17920 10198
rect 17868 10134 17920 10140
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17512 9722 17540 10066
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17512 9586 17540 9658
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 8974 17632 9318
rect 17880 8974 17908 9862
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17052 8634 17080 8910
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17604 8498 17632 8910
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17696 8566 17724 8774
rect 17880 8634 17908 8910
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17040 8492 17092 8498
rect 17224 8492 17276 8498
rect 17092 8452 17172 8480
rect 17040 8434 17092 8440
rect 17144 7750 17172 8452
rect 17224 8434 17276 8440
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17236 8401 17264 8434
rect 17222 8392 17278 8401
rect 17222 8327 17278 8336
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17144 6390 17172 7686
rect 17590 7576 17646 7585
rect 17590 7511 17646 7520
rect 17604 7410 17632 7511
rect 17696 7410 17724 7686
rect 17972 7546 18000 10678
rect 18144 10532 18196 10538
rect 18144 10474 18196 10480
rect 18156 10266 18184 10474
rect 18144 10260 18196 10266
rect 18144 10202 18196 10208
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 10062 18368 10202
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18432 9994 18460 10678
rect 18524 10538 18552 11086
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18524 10062 18552 10474
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18432 9722 18460 9930
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8634 18276 8774
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17972 7410 18000 7482
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17236 6866 17264 7142
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17512 6798 17540 7142
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17604 6730 17632 7346
rect 17788 7313 17816 7346
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17972 7002 18000 7346
rect 18064 7342 18092 7822
rect 18052 7336 18104 7342
rect 18696 7336 18748 7342
rect 18052 7278 18104 7284
rect 18510 7304 18566 7313
rect 18696 7278 18748 7284
rect 18510 7239 18566 7248
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17972 6866 18000 6938
rect 18524 6866 18552 7239
rect 18708 7002 18736 7278
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17236 6390 17264 6598
rect 17328 6458 17356 6598
rect 17604 6474 17632 6666
rect 17316 6452 17368 6458
rect 17604 6446 17724 6474
rect 17316 6394 17368 6400
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17144 6186 17172 6326
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16868 5766 16988 5794
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16868 5370 16896 5646
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16684 4622 16712 5170
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3398 16436 4014
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16592 3738 16620 3878
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16684 3670 16712 3878
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16684 3126 16712 3606
rect 16868 3466 16896 4558
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16500 2446 16528 2994
rect 16960 2774 16988 5766
rect 17052 5030 17080 6054
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17224 5704 17276 5710
rect 17224 5646 17276 5652
rect 17236 5234 17264 5646
rect 17328 5234 17356 5850
rect 17420 5710 17448 5850
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17408 5228 17460 5234
rect 17512 5216 17540 5578
rect 17604 5234 17632 6326
rect 17696 5710 17724 6446
rect 18248 6390 18276 6734
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5710 18276 6054
rect 18524 5914 18552 6802
rect 18616 6798 18644 6938
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18616 5302 18644 5782
rect 18604 5296 18656 5302
rect 18604 5238 18656 5244
rect 17460 5188 17540 5216
rect 17592 5228 17644 5234
rect 17408 5170 17460 5176
rect 18512 5228 18564 5234
rect 17644 5188 17724 5216
rect 17592 5170 17644 5176
rect 17236 5098 17264 5170
rect 17224 5092 17276 5098
rect 17224 5034 17276 5040
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4758 17172 4966
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17236 4282 17264 5034
rect 17328 4758 17356 5170
rect 17420 4826 17448 5170
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17328 4486 17356 4694
rect 17696 4554 17724 5188
rect 18512 5170 18564 5176
rect 18524 4826 18552 5170
rect 18800 5030 18828 18022
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18892 15706 18920 15914
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18892 14414 18920 15642
rect 18880 14408 18932 14414
rect 18880 14350 18932 14356
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18892 12442 18920 12718
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18878 10704 18934 10713
rect 18878 10639 18880 10648
rect 18932 10639 18934 10648
rect 18880 10610 18932 10616
rect 18892 10470 18920 10610
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18984 9382 19012 18142
rect 19260 17270 19288 19332
rect 19536 19360 19564 19751
rect 19628 19689 19656 19790
rect 19614 19680 19670 19689
rect 19614 19615 19670 19624
rect 19720 19378 19748 20420
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19812 19990 19840 20198
rect 19904 20058 19932 21898
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19996 20942 20024 21422
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19996 20602 20024 20878
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19892 20052 19944 20058
rect 19892 19994 19944 20000
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19904 19446 19932 19790
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19616 19372 19668 19378
rect 19536 19332 19616 19360
rect 19340 19314 19392 19320
rect 19616 19314 19668 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19996 18766 20024 20538
rect 20088 20346 20116 21966
rect 20180 21962 20208 22646
rect 20456 22574 20484 22918
rect 20640 22658 20668 24228
rect 21100 24138 21128 24278
rect 21284 24138 21312 24890
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20916 23730 20944 24006
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 20640 22642 20760 22658
rect 20640 22636 20772 22642
rect 20640 22630 20720 22636
rect 20720 22578 20772 22584
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20272 22030 20300 22510
rect 20536 22432 20588 22438
rect 20536 22374 20588 22380
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20548 22234 20576 22374
rect 20536 22228 20588 22234
rect 20536 22170 20588 22176
rect 20732 22166 20760 22374
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20168 20460 20220 20466
rect 20272 20448 20300 20742
rect 20220 20420 20300 20448
rect 20168 20402 20220 20408
rect 20088 20318 20208 20346
rect 20074 19952 20130 19961
rect 20180 19922 20208 20318
rect 20074 19887 20130 19896
rect 20168 19916 20220 19922
rect 20088 19854 20116 19887
rect 20168 19858 20220 19864
rect 20076 19848 20128 19854
rect 20180 19825 20208 19858
rect 20076 19790 20128 19796
rect 20166 19816 20222 19825
rect 20166 19751 20222 19760
rect 20364 19530 20392 21082
rect 20640 20874 20668 21830
rect 21008 21622 21036 22578
rect 21100 21690 21128 24074
rect 21376 23798 21404 24142
rect 21548 24064 21600 24070
rect 21548 24006 21600 24012
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21192 22778 21220 23666
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20812 21412 20864 21418
rect 20812 21354 20864 21360
rect 20824 20942 20852 21354
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20916 20806 20944 21490
rect 21100 21078 21128 21626
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20272 19502 20392 19530
rect 20456 19514 20484 19790
rect 20640 19514 20668 20402
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20444 19508 20496 19514
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 18834 20116 19314
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19248 17264 19300 17270
rect 19248 17206 19300 17212
rect 19352 16114 19380 18702
rect 20088 18426 20116 18770
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 20272 17746 20300 19502
rect 20444 19450 20496 19456
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20628 19372 20680 19378
rect 20732 19360 20760 20198
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 19378 20852 19654
rect 20680 19332 20760 19360
rect 20812 19372 20864 19378
rect 20628 19314 20680 19320
rect 20812 19314 20864 19320
rect 20364 18902 20392 19314
rect 20916 19258 20944 20742
rect 21008 19378 21036 20742
rect 21100 20466 21128 21014
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21192 20602 21220 20810
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21376 20466 21404 23734
rect 21560 23526 21588 24006
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21744 23322 21772 24754
rect 21824 24676 21876 24682
rect 21824 24618 21876 24624
rect 21836 24342 21864 24618
rect 22020 24342 22048 25230
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21836 23798 21864 24142
rect 21928 24070 21956 24142
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21824 23792 21876 23798
rect 21824 23734 21876 23740
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21744 23118 21772 23258
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21468 22642 21496 22918
rect 21744 22778 21772 23054
rect 22020 22982 22048 24278
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 21744 22642 21772 22714
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21744 22098 21772 22578
rect 21836 22098 21864 22918
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21744 21010 21772 22034
rect 22112 21690 22140 24210
rect 22100 21684 22152 21690
rect 22100 21626 22152 21632
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21192 19990 21220 20402
rect 21180 19984 21232 19990
rect 21180 19926 21232 19932
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 20824 19230 20944 19258
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19444 17134 19472 17682
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17338 19748 17478
rect 19996 17338 20024 17546
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19444 16046 19472 17070
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19248 16040 19300 16046
rect 19432 16040 19484 16046
rect 19248 15982 19300 15988
rect 19352 15988 19432 15994
rect 19352 15982 19484 15988
rect 19260 15162 19288 15982
rect 19352 15966 19472 15982
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19260 14940 19288 15098
rect 19352 15094 19380 15966
rect 19628 15910 19656 16186
rect 19720 16114 19748 16526
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19444 15502 19472 15846
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 19260 14912 19380 14940
rect 19352 13870 19380 14912
rect 19536 14550 19564 15438
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19444 14074 19472 14350
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19352 13326 19380 13806
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19444 13530 19472 13738
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19076 11150 19104 11698
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19076 10810 19104 11086
rect 19260 10810 19288 11698
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19444 10470 19472 13466
rect 19720 12986 19748 14350
rect 19812 13802 19840 17002
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 16114 20300 16594
rect 20352 16516 20404 16522
rect 20352 16458 20404 16464
rect 20364 16114 20392 16458
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20352 16108 20404 16114
rect 20352 16050 20404 16056
rect 20260 15972 20312 15978
rect 20260 15914 20312 15920
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19536 11354 19564 12038
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19720 10674 19748 12174
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19812 10810 19840 11018
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19432 10464 19484 10470
rect 19432 10406 19484 10412
rect 19340 10260 19392 10266
rect 19616 10260 19668 10266
rect 19392 10220 19616 10248
rect 19340 10202 19392 10208
rect 19616 10202 19668 10208
rect 19432 10124 19484 10130
rect 19260 10084 19432 10112
rect 19260 9518 19288 10084
rect 19432 10066 19484 10072
rect 19720 10062 19748 10610
rect 19904 10266 19932 15506
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19996 14074 20024 14282
rect 20088 14074 20116 14418
rect 20272 14278 20300 15914
rect 20364 15706 20392 16050
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20732 15502 20760 16186
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14272 20312 14278
rect 20260 14214 20312 14220
rect 20272 14074 20300 14214
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 19984 13796 20036 13802
rect 19984 13738 20036 13744
rect 19996 12306 20024 13738
rect 20456 13530 20484 14758
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20640 13326 20668 13942
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 20444 13252 20496 13258
rect 20444 13194 20496 13200
rect 20456 12850 20484 13194
rect 20640 12986 20668 13262
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 20364 12238 20392 12582
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20640 11778 20668 12922
rect 20732 12238 20760 13126
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20640 11762 20760 11778
rect 20640 11756 20772 11762
rect 20640 11750 20720 11756
rect 20720 11698 20772 11704
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11150 20024 11494
rect 20548 11354 20576 11630
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20548 11150 20576 11290
rect 20640 11150 20668 11630
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 19996 10742 20024 11086
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20180 10810 20208 10950
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20088 10266 20116 10542
rect 20180 10470 20208 10746
rect 20732 10742 20760 11698
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 19260 9110 19288 9454
rect 19248 9104 19300 9110
rect 19248 9046 19300 9052
rect 19260 8498 19288 9046
rect 20088 9024 20116 10202
rect 20272 9586 20300 10610
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20088 8996 20208 9024
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19720 8634 19748 8774
rect 20088 8634 20116 8842
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 7886 19288 8434
rect 20180 7954 20208 8996
rect 20272 8650 20300 9522
rect 20732 9042 20760 10678
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20272 8622 20392 8650
rect 20364 8498 20392 8622
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6474 19288 6734
rect 19352 6662 19380 7822
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19260 6446 19380 6474
rect 19352 6202 19380 6446
rect 19444 6322 19472 7686
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 19720 7410 19748 7482
rect 19904 7478 19932 7890
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19708 7404 19760 7410
rect 19760 7364 19840 7392
rect 19708 7346 19760 7352
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19536 6866 19564 7278
rect 19708 7200 19760 7206
rect 19628 7160 19708 7188
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19352 6174 19472 6202
rect 19248 5908 19300 5914
rect 19248 5850 19300 5856
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18984 5098 19012 5170
rect 19076 5098 19104 5646
rect 19260 5642 19288 5850
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19260 5216 19288 5578
rect 19340 5228 19392 5234
rect 19260 5188 19340 5216
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 19076 4622 19104 5034
rect 19260 4690 19288 5188
rect 19340 5170 19392 5176
rect 19444 4758 19472 6174
rect 19536 5710 19564 6802
rect 19628 6730 19656 7160
rect 19708 7142 19760 7148
rect 19812 6882 19840 7364
rect 19720 6866 19840 6882
rect 19708 6860 19840 6866
rect 19760 6854 19840 6860
rect 19708 6802 19760 6808
rect 19904 6798 19932 7414
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 6254 19748 6666
rect 19892 6316 19944 6322
rect 19996 6304 20024 7754
rect 20088 7546 20116 7822
rect 20168 7744 20220 7750
rect 20168 7686 20220 7692
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20074 7440 20130 7449
rect 20074 7375 20076 7384
rect 20128 7375 20130 7384
rect 20076 7346 20128 7352
rect 20088 6934 20116 7346
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20180 6662 20208 7686
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20272 6458 20300 8434
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20548 7886 20576 8230
rect 20640 7954 20668 8434
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20640 7546 20668 7890
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 19944 6276 20024 6304
rect 19892 6258 19944 6264
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19812 5914 19840 6190
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19904 5794 19932 6258
rect 20272 6186 20300 6394
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 19720 5766 19932 5794
rect 19982 5808 20038 5817
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5234 19564 5646
rect 19720 5574 19748 5766
rect 19982 5743 20038 5752
rect 19996 5710 20024 5743
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3398 17632 4082
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16592 2746 16988 2774
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 16132 800 16160 2382
rect 16592 2378 16620 2746
rect 17052 2650 17080 2994
rect 17604 2990 17632 3334
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17696 2582 17724 4490
rect 19076 4282 19104 4558
rect 19260 4282 19288 4626
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 17960 4004 18012 4010
rect 17960 3946 18012 3952
rect 17972 3738 18000 3946
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3738 18092 3878
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17880 3126 17908 3606
rect 18156 3466 18184 4082
rect 18248 3534 18276 4082
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 19338 3632 19394 3641
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 17868 3120 17920 3126
rect 18248 3074 18276 3470
rect 18432 3346 18460 3606
rect 19338 3567 19340 3576
rect 19392 3567 19394 3576
rect 19340 3538 19392 3544
rect 18604 3392 18656 3398
rect 18432 3340 18604 3346
rect 18432 3334 18656 3340
rect 18432 3318 18644 3334
rect 17868 3062 17920 3068
rect 18156 3046 18276 3074
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 18156 2990 18184 3046
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 17684 2576 17736 2582
rect 17684 2518 17736 2524
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 16580 2372 16632 2378
rect 16580 2314 16632 2320
rect 17420 800 17448 2382
rect 19352 2378 19380 3062
rect 19444 2990 19472 4558
rect 19432 2984 19484 2990
rect 19432 2926 19484 2932
rect 19444 2446 19472 2926
rect 19536 2650 19564 5170
rect 19720 4434 19748 5510
rect 20088 5234 20116 5510
rect 20180 5370 20208 6054
rect 20456 5710 20484 6258
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 19628 4406 19748 4434
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 18696 2372 18748 2378
rect 18696 2314 18748 2320
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 18708 800 18736 2314
rect 18880 2304 18932 2310
rect 18878 2272 18880 2281
rect 18932 2272 18934 2281
rect 18878 2207 18934 2216
rect 19628 1902 19656 4406
rect 20364 4282 20392 4558
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20456 4214 20484 4422
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19720 3670 19748 4014
rect 20732 3942 20760 8978
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 20732 3534 20760 3878
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20352 3460 20404 3466
rect 20352 3402 20404 3408
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19720 3126 19748 3334
rect 19708 3120 19760 3126
rect 19708 3062 19760 3068
rect 20364 2854 20392 3402
rect 20640 2990 20668 3402
rect 20732 3126 20760 3470
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 19616 1896 19668 1902
rect 19616 1838 19668 1844
rect 19996 800 20024 2382
rect 20824 2310 20852 19230
rect 21100 19174 21128 19790
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18970 21128 19110
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20916 16114 20944 16730
rect 21008 16590 21036 18362
rect 21192 18290 21220 19926
rect 21376 19854 21404 20402
rect 21744 20058 21772 20810
rect 21836 20398 21864 21490
rect 22112 21162 22140 21626
rect 22112 21134 22324 21162
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 21824 20392 21876 20398
rect 21824 20334 21876 20340
rect 22112 20380 22140 20946
rect 22192 20392 22244 20398
rect 22112 20352 22192 20380
rect 21732 20052 21784 20058
rect 21732 19994 21784 20000
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21928 19854 21956 19926
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21376 19446 21404 19790
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21824 19712 21876 19718
rect 21824 19654 21876 19660
rect 21652 19514 21680 19654
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21376 18426 21404 18702
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21192 16658 21220 18226
rect 21284 17542 21312 18226
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 16794 21312 17478
rect 21376 17338 21404 18362
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21364 17196 21416 17202
rect 21364 17138 21416 17144
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 21376 16658 21404 17138
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20916 15162 20944 16050
rect 21192 16046 21220 16594
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21468 16402 21496 19314
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 21560 17338 21588 18226
rect 21652 18154 21680 18770
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 21836 17678 21864 19654
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 21928 17882 21956 18226
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21652 17202 21680 17614
rect 21732 17264 21784 17270
rect 21732 17206 21784 17212
rect 21640 17196 21692 17202
rect 21560 17156 21640 17184
rect 21560 16522 21588 17156
rect 21640 17138 21692 17144
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21652 16590 21680 16934
rect 21640 16584 21692 16590
rect 21744 16572 21772 17206
rect 21916 17196 21968 17202
rect 22020 17184 22048 18022
rect 22112 17746 22140 20352
rect 22192 20334 22244 20340
rect 22296 19922 22324 21134
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22204 18154 22232 18702
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 22112 17338 22140 17478
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22388 17252 22416 30058
rect 23940 30048 23992 30054
rect 23940 29990 23992 29996
rect 24124 30048 24176 30054
rect 24124 29990 24176 29996
rect 26148 30048 26200 30054
rect 26148 29990 26200 29996
rect 23480 29028 23532 29034
rect 23480 28970 23532 28976
rect 23492 28490 23520 28970
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23480 28076 23532 28082
rect 23480 28018 23532 28024
rect 23492 27538 23520 28018
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22572 27130 22600 27338
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 23492 26926 23520 27474
rect 23480 26920 23532 26926
rect 23400 26868 23480 26874
rect 23400 26862 23532 26868
rect 23400 26846 23520 26862
rect 23296 26512 23348 26518
rect 23296 26454 23348 26460
rect 23308 25974 23336 26454
rect 23400 26382 23428 26846
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23492 26314 23520 26726
rect 23676 26314 23704 27950
rect 23848 27872 23900 27878
rect 23848 27814 23900 27820
rect 23860 27674 23888 27814
rect 23848 27668 23900 27674
rect 23848 27610 23900 27616
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23768 26586 23796 26862
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23952 26330 23980 29990
rect 24032 28552 24084 28558
rect 24032 28494 24084 28500
rect 24044 28014 24072 28494
rect 24032 28008 24084 28014
rect 24032 27950 24084 27956
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23664 26308 23716 26314
rect 23952 26302 24072 26330
rect 23664 26250 23716 26256
rect 23940 26240 23992 26246
rect 23768 26200 23940 26228
rect 23296 25968 23348 25974
rect 23296 25910 23348 25916
rect 23768 25294 23796 26200
rect 23940 26182 23992 26188
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23756 25288 23808 25294
rect 24044 25242 24072 26302
rect 23756 25230 23808 25236
rect 23112 25152 23164 25158
rect 23112 25094 23164 25100
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22572 24410 22600 24822
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22848 24410 22876 24686
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 23124 24342 23152 25094
rect 23584 24750 23612 25230
rect 23768 24886 23796 25230
rect 23860 25214 24072 25242
rect 23756 24880 23808 24886
rect 23756 24822 23808 24828
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23112 24336 23164 24342
rect 23112 24278 23164 24284
rect 23676 24138 23704 24550
rect 23768 24274 23796 24822
rect 23756 24268 23808 24274
rect 23756 24210 23808 24216
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 23860 23254 23888 25214
rect 24032 25152 24084 25158
rect 24032 25094 24084 25100
rect 24044 24886 24072 25094
rect 24032 24880 24084 24886
rect 24032 24822 24084 24828
rect 24044 24206 24072 24822
rect 24032 24200 24084 24206
rect 24032 24142 24084 24148
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23848 23248 23900 23254
rect 23848 23190 23900 23196
rect 23572 23180 23624 23186
rect 23572 23122 23624 23128
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23400 22166 23428 22714
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22480 20602 22508 20810
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22572 20466 22600 22034
rect 23584 21962 23612 23122
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 22940 21554 22968 21830
rect 23124 21554 23152 21830
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23204 21548 23256 21554
rect 23204 21490 23256 21496
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23124 20874 23152 21490
rect 23216 21146 23244 21490
rect 23204 21140 23256 21146
rect 23204 21082 23256 21088
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23492 20806 23520 21490
rect 23584 21078 23612 21898
rect 23676 21554 23704 22986
rect 23860 22234 23888 23190
rect 23952 22710 23980 24074
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23848 22228 23900 22234
rect 23848 22170 23900 22176
rect 23860 22094 23888 22170
rect 23860 22066 23980 22094
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23572 21072 23624 21078
rect 23572 21014 23624 21020
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22572 20330 22600 20402
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22848 19514 22876 19790
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22480 18970 22508 19246
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22848 18766 22876 19450
rect 23308 19446 23336 19858
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 23308 18290 23336 19382
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 22204 17224 22416 17252
rect 21968 17156 22048 17184
rect 22100 17196 22152 17202
rect 21916 17138 21968 17144
rect 22100 17138 22152 17144
rect 21824 16584 21876 16590
rect 21744 16544 21824 16572
rect 21640 16526 21692 16532
rect 21824 16526 21876 16532
rect 21548 16516 21600 16522
rect 21548 16458 21600 16464
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21284 15706 21312 16390
rect 21468 16374 21588 16402
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20916 14958 20944 15098
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21008 14074 21036 14282
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20916 12986 20944 13194
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 21008 12850 21036 13874
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21284 11694 21312 12854
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 20904 11280 20956 11286
rect 21560 11234 21588 16374
rect 21928 15978 21956 17138
rect 22112 16454 22140 17138
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22008 16040 22060 16046
rect 22008 15982 22060 15988
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 22020 15434 22048 15982
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22020 15026 22048 15370
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22112 14822 22140 15846
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22008 13864 22060 13870
rect 22060 13824 22140 13852
rect 22008 13806 22060 13812
rect 22112 13734 22140 13824
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 22008 13456 22060 13462
rect 22008 13398 22060 13404
rect 21916 13252 21968 13258
rect 21916 13194 21968 13200
rect 21928 12986 21956 13194
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 12850 22048 13398
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22112 12782 22140 13670
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 21640 12232 21692 12238
rect 22008 12232 22060 12238
rect 21640 12174 21692 12180
rect 21836 12192 22008 12220
rect 20904 11222 20956 11228
rect 20916 9722 20944 11222
rect 21376 11206 21588 11234
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21284 10810 21312 11018
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 21192 9586 21220 10610
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 21100 8974 21128 9386
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20916 8294 20944 8774
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 20916 7478 20944 8230
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 20904 7472 20956 7478
rect 20904 7414 20956 7420
rect 21008 7410 21036 7890
rect 21284 7886 21312 8026
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 21008 5574 21036 7346
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 5710 21128 6598
rect 21192 6254 21220 7142
rect 21376 6662 21404 11206
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21560 10810 21588 11086
rect 21652 11082 21680 12174
rect 21836 11558 21864 12192
rect 22008 12174 22060 12180
rect 21916 11620 21968 11626
rect 21916 11562 21968 11568
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21732 11280 21784 11286
rect 21732 11222 21784 11228
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21652 10674 21680 11018
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21560 9586 21588 10474
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21652 9722 21680 10066
rect 21744 10062 21772 11222
rect 21836 11082 21864 11494
rect 21928 11286 21956 11562
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21824 11076 21876 11082
rect 21824 11018 21876 11024
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21640 9716 21692 9722
rect 21640 9658 21692 9664
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21836 8022 21864 11018
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21928 8294 21956 9454
rect 22112 9330 22140 9590
rect 22020 9302 22140 9330
rect 22020 9178 22048 9302
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21468 7410 21496 7754
rect 21560 7478 21588 7754
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21836 7410 21864 7958
rect 22112 7886 22140 9114
rect 22204 9110 22232 17224
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16658 22416 16934
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22480 16250 22508 16526
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22296 14958 22324 15574
rect 22388 15502 22416 16050
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22468 15360 22520 15366
rect 23204 15360 23256 15366
rect 22520 15320 22600 15348
rect 22468 15302 22520 15308
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 13802 22324 14214
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22388 12918 22416 13126
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22296 11218 22324 12174
rect 22388 11558 22416 12854
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22388 10606 22416 11494
rect 22480 11218 22508 12174
rect 22572 11354 22600 15320
rect 23204 15302 23256 15308
rect 23216 15094 23244 15302
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 22928 14884 22980 14890
rect 22928 14826 22980 14832
rect 22940 14074 22968 14826
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23480 14000 23532 14006
rect 23480 13942 23532 13948
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23216 12238 23244 13806
rect 23492 13530 23520 13942
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23584 12764 23612 15506
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 15162 23704 15438
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23664 12776 23716 12782
rect 23584 12736 23664 12764
rect 23664 12718 23716 12724
rect 23676 12306 23704 12718
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22848 11218 22876 12174
rect 23480 11620 23532 11626
rect 23480 11562 23532 11568
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 11354 23060 11494
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 23492 11218 23520 11562
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22204 8566 22232 9046
rect 22388 8974 22416 10542
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22296 7886 22324 8026
rect 22388 7886 22416 8910
rect 22848 8090 22876 11154
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 23216 10606 23244 11018
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23124 10266 23152 10542
rect 23112 10260 23164 10266
rect 23112 10202 23164 10208
rect 23216 10130 23244 10542
rect 23676 10130 23704 12242
rect 23204 10124 23256 10130
rect 23124 10084 23204 10112
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22652 8016 22704 8022
rect 22704 7976 22784 8004
rect 22652 7958 22704 7964
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22100 7880 22152 7886
rect 22284 7880 22336 7886
rect 22100 7822 22152 7828
rect 22204 7828 22284 7834
rect 22204 7822 22336 7828
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22204 7806 22324 7822
rect 22572 7818 22600 7890
rect 22756 7886 22784 7976
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22560 7812 22612 7818
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22112 7546 22140 7686
rect 22100 7540 22152 7546
rect 22100 7482 22152 7488
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21640 6384 21692 6390
rect 21640 6326 21692 6332
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 21100 3942 21128 4966
rect 21192 4554 21220 6190
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21272 5568 21324 5574
rect 21272 5510 21324 5516
rect 21284 5234 21312 5510
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21376 5030 21404 5646
rect 21468 5642 21496 6258
rect 21560 5846 21588 6258
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21652 5574 21680 6326
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21836 5778 21864 6258
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21928 4690 21956 7414
rect 22204 5370 22232 7806
rect 22560 7754 22612 7760
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 7546 22324 7686
rect 22664 7546 22692 7822
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22848 7410 22876 8026
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22940 7290 22968 9590
rect 23124 9042 23152 10084
rect 23204 10066 23256 10072
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23768 9654 23796 21286
rect 23952 21010 23980 22066
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 24044 16182 24072 16390
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 24136 12434 24164 29990
rect 25320 28688 25372 28694
rect 25320 28630 25372 28636
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24228 28082 24256 28358
rect 24504 28218 24532 28494
rect 24492 28212 24544 28218
rect 24492 28154 24544 28160
rect 25136 28144 25188 28150
rect 25136 28086 25188 28092
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24768 28008 24820 28014
rect 24768 27950 24820 27956
rect 25044 28008 25096 28014
rect 25044 27950 25096 27956
rect 24780 27470 24808 27950
rect 25056 27674 25084 27950
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25148 27470 25176 28086
rect 25332 27470 25360 28630
rect 25504 28552 25556 28558
rect 25504 28494 25556 28500
rect 25516 27878 25544 28494
rect 25780 28484 25832 28490
rect 25780 28426 25832 28432
rect 25792 28014 25820 28426
rect 25964 28416 26016 28422
rect 25964 28358 26016 28364
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25504 27872 25556 27878
rect 25504 27814 25556 27820
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 25320 27464 25372 27470
rect 25320 27406 25372 27412
rect 24492 27056 24544 27062
rect 24492 26998 24544 27004
rect 24504 26042 24532 26998
rect 24780 26790 24808 27406
rect 25516 27402 25544 27814
rect 25792 27674 25820 27950
rect 25780 27668 25832 27674
rect 25780 27610 25832 27616
rect 25976 27402 26004 28358
rect 25504 27396 25556 27402
rect 25504 27338 25556 27344
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24780 26450 24808 26726
rect 24964 26586 24992 26862
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 25884 26450 25912 27338
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 25872 26444 25924 26450
rect 25872 26386 25924 26392
rect 24492 26036 24544 26042
rect 24492 25978 24544 25984
rect 24780 25906 24808 26386
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 25240 26042 25268 26250
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25884 25974 25912 26386
rect 25872 25968 25924 25974
rect 25872 25910 25924 25916
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 24228 24410 24256 24686
rect 25148 24410 25176 24822
rect 24216 24404 24268 24410
rect 24216 24346 24268 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25688 24132 25740 24138
rect 25688 24074 25740 24080
rect 25700 23866 25728 24074
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25228 23792 25280 23798
rect 25228 23734 25280 23740
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 25056 22642 25084 22918
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24228 13258 24256 21490
rect 24412 20942 24440 22374
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 24504 21690 24532 22034
rect 25240 22001 25268 23734
rect 25412 23044 25464 23050
rect 25412 22986 25464 22992
rect 25424 22778 25452 22986
rect 25412 22772 25464 22778
rect 25412 22714 25464 22720
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 25226 21992 25282 22001
rect 25226 21927 25282 21936
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 26068 21418 26096 22034
rect 26056 21412 26108 21418
rect 26056 21354 26108 21360
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24504 20602 24532 20878
rect 25332 20874 25360 21286
rect 25320 20868 25372 20874
rect 25320 20810 25372 20816
rect 26068 20806 26096 21354
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 26056 20800 26108 20806
rect 26056 20742 26108 20748
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24596 17882 24624 18294
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24688 17678 24716 19314
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24504 16182 24532 16662
rect 24688 16590 24716 17614
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 24688 16250 24716 16526
rect 24676 16244 24728 16250
rect 24676 16186 24728 16192
rect 24492 16176 24544 16182
rect 24492 16118 24544 16124
rect 24688 15502 24716 16186
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24400 15360 24452 15366
rect 24400 15302 24452 15308
rect 24412 15026 24440 15302
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24216 13252 24268 13258
rect 24216 13194 24268 13200
rect 24044 12406 24164 12434
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23952 11694 23980 12038
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23756 9648 23808 9654
rect 23756 9590 23808 9596
rect 23572 9580 23624 9586
rect 23572 9522 23624 9528
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23112 9036 23164 9042
rect 23112 8978 23164 8984
rect 23400 8974 23428 9318
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23308 8430 23336 8842
rect 23492 8634 23520 8910
rect 23584 8838 23612 9522
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23584 8514 23612 8774
rect 23676 8634 23704 9454
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23584 8498 23704 8514
rect 23480 8492 23532 8498
rect 23584 8492 23716 8498
rect 23584 8486 23664 8492
rect 23480 8434 23532 8440
rect 23664 8434 23716 8440
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23204 7880 23256 7886
rect 23308 7834 23336 8366
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23400 7886 23428 8230
rect 23492 7970 23520 8434
rect 23860 8362 23888 8842
rect 24044 8650 24072 12406
rect 24228 11830 24256 13194
rect 24492 12096 24544 12102
rect 24492 12038 24544 12044
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24504 11558 24532 12038
rect 24492 11552 24544 11558
rect 24492 11494 24544 11500
rect 24504 11218 24532 11494
rect 24492 11212 24544 11218
rect 24492 11154 24544 11160
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 24136 10266 24164 10678
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24216 9648 24268 9654
rect 24216 9590 24268 9596
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 23952 8622 24072 8650
rect 24136 8634 24164 9522
rect 24124 8628 24176 8634
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23860 7970 23888 8298
rect 23492 7942 23612 7970
rect 23256 7828 23336 7834
rect 23204 7822 23336 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23216 7806 23336 7822
rect 23308 7410 23336 7806
rect 23492 7449 23520 7822
rect 23478 7440 23534 7449
rect 23296 7404 23348 7410
rect 23478 7375 23534 7384
rect 23296 7346 23348 7352
rect 22848 7262 22968 7290
rect 23112 7336 23164 7342
rect 23584 7290 23612 7942
rect 23112 7278 23164 7284
rect 22848 6322 22876 7262
rect 22560 6316 22612 6322
rect 22560 6258 22612 6264
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22572 5914 22600 6258
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3602 21128 3878
rect 21088 3596 21140 3602
rect 21088 3538 21140 3544
rect 21192 2582 21220 4490
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21284 3194 21312 3402
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 21928 1970 21956 4626
rect 22296 3670 22324 5170
rect 22480 4758 22508 5170
rect 22664 4758 22692 5170
rect 22756 4826 22784 5170
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22468 4752 22520 4758
rect 22468 4694 22520 4700
rect 22652 4752 22704 4758
rect 22652 4694 22704 4700
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22572 3670 22600 3878
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22468 3664 22520 3670
rect 22468 3606 22520 3612
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 22480 3534 22508 3606
rect 22468 3528 22520 3534
rect 22664 3482 22692 3878
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22468 3470 22520 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 3194 22048 3402
rect 22480 3398 22508 3470
rect 22572 3454 22692 3482
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22572 3058 22600 3454
rect 22756 3058 22784 3538
rect 22848 3398 22876 4558
rect 22940 3942 22968 5646
rect 23124 4622 23152 7278
rect 23492 7262 23612 7290
rect 23768 7942 23888 7970
rect 23492 6338 23520 7262
rect 23216 6322 23520 6338
rect 23768 6322 23796 7942
rect 23848 7812 23900 7818
rect 23848 7754 23900 7760
rect 23860 7342 23888 7754
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23952 6730 23980 8622
rect 24124 8570 24176 8576
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 24044 8090 24072 8434
rect 24124 8356 24176 8362
rect 24124 8298 24176 8304
rect 24136 8090 24164 8298
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 24228 7970 24256 9590
rect 24504 8974 24532 11154
rect 24872 9382 24900 20742
rect 24952 20392 25004 20398
rect 24952 20334 25004 20340
rect 24964 19378 24992 20334
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 25148 19514 25176 19722
rect 25976 19514 26004 19722
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 26068 19310 26096 20742
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 16454 25084 18158
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 17610 25544 18022
rect 25504 17604 25556 17610
rect 25504 17546 25556 17552
rect 25596 17196 25648 17202
rect 25596 17138 25648 17144
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25044 16448 25096 16454
rect 25044 16390 25096 16396
rect 25056 16114 25084 16390
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25148 16046 25176 16594
rect 25424 16114 25452 16934
rect 25608 16794 25636 17138
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 26068 16658 26096 17070
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25516 16250 25544 16458
rect 26068 16454 26096 16594
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 25148 14958 25176 15982
rect 26068 14958 26096 16390
rect 25136 14952 25188 14958
rect 25136 14894 25188 14900
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25148 14482 25176 14894
rect 25412 14816 25464 14822
rect 25412 14758 25464 14764
rect 25136 14476 25188 14482
rect 25136 14418 25188 14424
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24964 12986 24992 13806
rect 25148 13734 25176 14418
rect 25424 14346 25452 14758
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25148 13394 25176 13670
rect 26068 13530 26096 13874
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25148 12238 25176 13330
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 12306 25728 12582
rect 26160 12434 26188 29990
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 26042 26280 26250
rect 26240 26036 26292 26042
rect 26240 25978 26292 25984
rect 26240 25900 26292 25906
rect 26240 25842 26292 25848
rect 26252 25226 26280 25842
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 26252 24818 26280 25162
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26252 23118 26280 24346
rect 26344 24138 26372 24550
rect 26332 24132 26384 24138
rect 26332 24074 26384 24080
rect 26528 24070 26556 30126
rect 27804 30116 27856 30122
rect 27804 30058 27856 30064
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 27080 27470 27108 28494
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27160 28416 27212 28422
rect 27160 28358 27212 28364
rect 27172 28082 27200 28358
rect 27160 28076 27212 28082
rect 27160 28018 27212 28024
rect 27356 28014 27384 28426
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27068 27464 27120 27470
rect 27068 27406 27120 27412
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27080 26994 27108 27406
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 26976 26376 27028 26382
rect 27344 26376 27396 26382
rect 26976 26318 27028 26324
rect 27172 26324 27344 26330
rect 27172 26318 27396 26324
rect 26792 26240 26844 26246
rect 26988 26228 27016 26318
rect 27172 26302 27384 26318
rect 27172 26228 27200 26302
rect 26988 26200 27200 26228
rect 26792 26182 26844 26188
rect 26804 25770 26832 26182
rect 27172 25906 27200 26200
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 27356 25974 27384 26182
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 26792 25764 26844 25770
rect 26792 25706 26844 25712
rect 27172 25294 27200 25842
rect 27356 25294 27384 25910
rect 27448 25498 27476 26862
rect 27632 25838 27660 27406
rect 27816 26330 27844 30058
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 27896 27396 27948 27402
rect 27896 27338 27948 27344
rect 27908 27130 27936 27338
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 27896 27124 27948 27130
rect 27896 27066 27948 27072
rect 28000 26994 28028 27270
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 28000 26518 28028 26930
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 27816 26302 27936 26330
rect 27804 26240 27856 26246
rect 27804 26182 27856 26188
rect 27816 26042 27844 26182
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 27620 25832 27672 25838
rect 27620 25774 27672 25780
rect 27436 25492 27488 25498
rect 27436 25434 27488 25440
rect 26792 25288 26844 25294
rect 26792 25230 26844 25236
rect 27160 25288 27212 25294
rect 27160 25230 27212 25236
rect 27344 25288 27396 25294
rect 27344 25230 27396 25236
rect 26804 24614 26832 25230
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 26792 24608 26844 24614
rect 26792 24550 26844 24556
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26804 23730 26832 24550
rect 27172 23730 27200 24754
rect 27448 24410 27476 24754
rect 27436 24404 27488 24410
rect 27436 24346 27488 24352
rect 27448 23730 27476 24346
rect 27540 24070 27568 24822
rect 27632 24818 27660 25774
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 27724 25294 27752 25638
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27620 24812 27672 24818
rect 27620 24754 27672 24760
rect 27632 24206 27660 24754
rect 27804 24676 27856 24682
rect 27804 24618 27856 24624
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27540 23730 27568 24006
rect 26792 23724 26844 23730
rect 26792 23666 26844 23672
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27528 23724 27580 23730
rect 27528 23666 27580 23672
rect 27172 23118 27200 23666
rect 27344 23656 27396 23662
rect 27344 23598 27396 23604
rect 27356 23118 27384 23598
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 27160 23112 27212 23118
rect 27160 23054 27212 23060
rect 27344 23112 27396 23118
rect 27344 23054 27396 23060
rect 26252 22642 26280 23054
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26700 22432 26752 22438
rect 26700 22374 26752 22380
rect 26608 22024 26660 22030
rect 26528 21984 26608 22012
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26252 21554 26280 21626
rect 26332 21616 26384 21622
rect 26332 21558 26384 21564
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 26344 21010 26372 21558
rect 26424 21548 26476 21554
rect 26528 21536 26556 21984
rect 26608 21966 26660 21972
rect 26712 21962 26740 22374
rect 27172 22234 27200 23054
rect 27632 22574 27660 24142
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27724 23322 27752 23598
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 27816 23202 27844 24618
rect 27908 23526 27936 26302
rect 27988 25832 28040 25838
rect 27988 25774 28040 25780
rect 28000 25498 28028 25774
rect 27988 25492 28040 25498
rect 27988 25434 28040 25440
rect 27896 23520 27948 23526
rect 27896 23462 27948 23468
rect 27724 23174 27844 23202
rect 27724 23050 27752 23174
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27724 22778 27752 22986
rect 27896 22976 27948 22982
rect 27896 22918 27948 22924
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 27908 22710 27936 22918
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27172 22094 27200 22170
rect 26988 22066 27200 22094
rect 26700 21956 26752 21962
rect 26700 21898 26752 21904
rect 26988 21554 27016 22066
rect 27068 21888 27120 21894
rect 27068 21830 27120 21836
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 26476 21508 26556 21536
rect 26976 21548 27028 21554
rect 26424 21490 26476 21496
rect 26976 21490 27028 21496
rect 26436 21146 26464 21490
rect 26424 21140 26476 21146
rect 26424 21082 26476 21088
rect 26332 21004 26384 21010
rect 26252 20964 26332 20992
rect 26252 19922 26280 20964
rect 26332 20946 26384 20952
rect 27080 20942 27108 21830
rect 27172 21690 27200 21830
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 27172 20874 27200 21626
rect 27528 21548 27580 21554
rect 27632 21536 27660 22510
rect 27580 21508 27660 21536
rect 27528 21490 27580 21496
rect 27344 21412 27396 21418
rect 27344 21354 27396 21360
rect 27356 21146 27384 21354
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 27160 20868 27212 20874
rect 27160 20810 27212 20816
rect 26344 20602 26372 20810
rect 26332 20596 26384 20602
rect 26332 20538 26384 20544
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27540 20058 27568 20402
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27632 19922 27660 21508
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26252 18290 26280 19314
rect 26804 19242 26832 19654
rect 26896 19242 26924 19858
rect 26976 19848 27028 19854
rect 27028 19808 27200 19836
rect 26976 19790 27028 19796
rect 27172 19378 27200 19808
rect 27252 19780 27304 19786
rect 27252 19722 27304 19728
rect 27264 19514 27292 19722
rect 27356 19514 27384 19858
rect 27252 19508 27304 19514
rect 27252 19450 27304 19456
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26884 19236 26936 19242
rect 26884 19178 26936 19184
rect 27172 18698 27200 19314
rect 27528 19236 27580 19242
rect 27528 19178 27580 19184
rect 27540 18698 27568 19178
rect 26792 18692 26844 18698
rect 26792 18634 26844 18640
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26332 18216 26384 18222
rect 26332 18158 26384 18164
rect 26240 18080 26292 18086
rect 26240 18022 26292 18028
rect 26252 17610 26280 18022
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 26344 17542 26372 18158
rect 26804 17610 26832 18634
rect 27540 18426 27568 18634
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27632 18290 27660 19858
rect 27724 19514 27752 20334
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27908 19922 27936 20198
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27724 18748 27752 19450
rect 27804 18760 27856 18766
rect 27724 18720 27804 18748
rect 27804 18702 27856 18708
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 27908 18358 27936 18566
rect 27896 18352 27948 18358
rect 27896 18294 27948 18300
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27436 17808 27488 17814
rect 27436 17750 27488 17756
rect 26792 17604 26844 17610
rect 26792 17546 26844 17552
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17202 26372 17478
rect 26804 17270 26832 17546
rect 27160 17536 27212 17542
rect 27160 17478 27212 17484
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 26792 17264 26844 17270
rect 26792 17206 26844 17212
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 27080 16658 27108 17274
rect 27172 16658 27200 17478
rect 27448 16794 27476 17750
rect 27632 17746 27660 18226
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27540 16674 27568 17614
rect 27632 17270 27660 17682
rect 27712 17536 27764 17542
rect 27712 17478 27764 17484
rect 27724 17270 27752 17478
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27448 16658 27568 16674
rect 27068 16652 27120 16658
rect 27068 16594 27120 16600
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 27436 16652 27568 16658
rect 27488 16646 27568 16652
rect 27436 16594 27488 16600
rect 26424 16516 26476 16522
rect 26424 16458 26476 16464
rect 26436 16250 26464 16458
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 27448 16182 27476 16594
rect 27896 16244 27948 16250
rect 27896 16186 27948 16192
rect 27436 16176 27488 16182
rect 27436 16118 27488 16124
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26252 15026 26280 16050
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27620 16040 27672 16046
rect 27620 15982 27672 15988
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 26240 15020 26292 15026
rect 26292 14980 26372 15008
rect 26240 14962 26292 14968
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26252 14414 26280 14758
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26344 13326 26372 14980
rect 27172 14958 27200 15370
rect 27264 15366 27292 15982
rect 27344 15496 27396 15502
rect 27344 15438 27396 15444
rect 27252 15360 27304 15366
rect 27252 15302 27304 15308
rect 27356 14958 27384 15438
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27436 14952 27488 14958
rect 27436 14894 27488 14900
rect 27172 14346 27200 14894
rect 27356 14346 27384 14894
rect 27448 14618 27476 14894
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27632 14414 27660 15982
rect 27908 15162 27936 16186
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27988 15156 28040 15162
rect 27988 15098 28040 15104
rect 28000 14906 28028 15098
rect 27724 14878 28028 14906
rect 27724 14618 27752 14878
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27172 13870 27200 14282
rect 27160 13864 27212 13870
rect 27160 13806 27212 13812
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26332 13320 26384 13326
rect 26332 13262 26384 13268
rect 26436 12986 26464 13670
rect 27172 13530 27200 13806
rect 27528 13796 27580 13802
rect 27528 13738 27580 13744
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 27160 13320 27212 13326
rect 27160 13262 27212 13268
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26620 12850 26648 13126
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26068 12406 26188 12434
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 25136 12232 25188 12238
rect 25136 12174 25188 12180
rect 25148 11642 25176 12174
rect 25056 11614 25176 11642
rect 25056 10606 25084 11614
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10742 25360 10950
rect 25320 10736 25372 10742
rect 25320 10678 25372 10684
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25056 9518 25084 10542
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24676 8832 24728 8838
rect 24676 8774 24728 8780
rect 24044 7942 24256 7970
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 23204 6316 23532 6322
rect 23256 6310 23480 6316
rect 23204 6258 23256 6264
rect 23480 6258 23532 6264
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 23768 5778 23796 6258
rect 23756 5772 23808 5778
rect 23756 5714 23808 5720
rect 23860 5710 23888 6258
rect 23940 6180 23992 6186
rect 23940 6122 23992 6128
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23952 5370 23980 6122
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 23848 5228 23900 5234
rect 23848 5170 23900 5176
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23480 4616 23532 4622
rect 23664 4616 23716 4622
rect 23532 4564 23664 4570
rect 23480 4558 23716 4564
rect 23124 4162 23152 4558
rect 23492 4542 23704 4558
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23032 4134 23152 4162
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3176 22876 3334
rect 22928 3188 22980 3194
rect 22848 3148 22928 3176
rect 22928 3130 22980 3136
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 22928 2916 22980 2922
rect 22928 2858 22980 2864
rect 22020 2825 22048 2858
rect 22006 2816 22062 2825
rect 22006 2751 22062 2760
rect 22940 2530 22968 2858
rect 23032 2774 23060 4134
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23124 3641 23152 3674
rect 23110 3632 23166 3641
rect 23110 3567 23166 3576
rect 23032 2746 23152 2774
rect 23124 2650 23152 2746
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23216 2530 23244 4422
rect 23768 4214 23796 4422
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23296 4072 23348 4078
rect 23860 4026 23888 5170
rect 23296 4014 23348 4020
rect 23308 3058 23336 4014
rect 23768 3998 23888 4026
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23400 3738 23428 3878
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23388 3596 23440 3602
rect 23388 3538 23440 3544
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23400 2938 23428 3538
rect 23676 3534 23704 3674
rect 23768 3534 23796 3998
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23492 3126 23520 3334
rect 23768 3194 23796 3470
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23308 2910 23428 2938
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23308 2650 23336 2910
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 22940 2502 23244 2530
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 22572 800 22600 2382
rect 23124 2378 23152 2502
rect 23296 2440 23348 2446
rect 23216 2400 23296 2428
rect 23112 2372 23164 2378
rect 23112 2314 23164 2320
rect 23216 800 23244 2400
rect 23296 2382 23348 2388
rect 23400 2378 23428 2790
rect 23584 2650 23612 2926
rect 24044 2825 24072 7942
rect 24688 7886 24716 8774
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 24964 7886 24992 8570
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24676 7880 24728 7886
rect 24676 7822 24728 7828
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24228 7546 24256 7822
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24320 6322 24348 7754
rect 24412 7410 24440 7822
rect 24688 7478 24716 7822
rect 24676 7472 24728 7478
rect 24676 7414 24728 7420
rect 24400 7404 24452 7410
rect 24452 7364 24532 7392
rect 24400 7346 24452 7352
rect 24504 6458 24532 7364
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24492 6452 24544 6458
rect 24492 6394 24544 6400
rect 24504 6322 24532 6394
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24136 4826 24164 6258
rect 24596 6186 24624 7278
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 24596 5710 24624 6122
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24780 5710 24808 6054
rect 24964 5710 24992 6054
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24124 4616 24176 4622
rect 24124 4558 24176 4564
rect 24136 4078 24164 4558
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24504 4214 24532 4422
rect 24492 4208 24544 4214
rect 24492 4150 24544 4156
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24136 3534 24164 4014
rect 25056 3942 25084 9454
rect 26068 7993 26096 12406
rect 26896 12220 26924 13262
rect 27068 13252 27120 13258
rect 27068 13194 27120 13200
rect 27080 12850 27108 13194
rect 27172 12986 27200 13262
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27172 12850 27200 12922
rect 27264 12850 27292 13126
rect 27540 12986 27568 13738
rect 27632 13462 27660 14350
rect 27896 13728 27948 13734
rect 27896 13670 27948 13676
rect 27620 13456 27672 13462
rect 27620 13398 27672 13404
rect 27632 13326 27660 13398
rect 27908 13394 27936 13670
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27448 12442 27476 12786
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 26976 12232 27028 12238
rect 26896 12192 26976 12220
rect 26896 11762 26924 12192
rect 26976 12174 27028 12180
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26884 11756 26936 11762
rect 26884 11698 26936 11704
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 26436 11150 26464 11698
rect 27540 11354 27568 11698
rect 27632 11694 27660 13262
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27724 12782 27752 13126
rect 27988 12844 28040 12850
rect 27988 12786 28040 12792
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 28000 11898 28028 12786
rect 28092 12434 28120 29990
rect 28552 29646 28580 31311
rect 28906 30016 28962 30025
rect 28906 29951 28962 29960
rect 28920 29646 28948 29951
rect 29012 29646 29040 32247
rect 29380 30258 29408 32671
rect 30286 32247 30342 33047
rect 30300 30326 30328 32247
rect 30288 30320 30340 30326
rect 30288 30262 30340 30268
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29736 30184 29788 30190
rect 29736 30126 29788 30132
rect 28540 29640 28592 29646
rect 28540 29582 28592 29588
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 28356 29572 28408 29578
rect 28356 29514 28408 29520
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28184 23866 28212 24074
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28172 23180 28224 23186
rect 28172 23122 28224 23128
rect 28184 16590 28212 23122
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28172 14884 28224 14890
rect 28172 14826 28224 14832
rect 28184 14346 28212 14826
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 28276 14618 28304 14758
rect 28264 14612 28316 14618
rect 28264 14554 28316 14560
rect 28172 14340 28224 14346
rect 28172 14282 28224 14288
rect 28092 12406 28212 12434
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 26148 11144 26200 11150
rect 26424 11144 26476 11150
rect 26200 11092 26280 11098
rect 26148 11086 26280 11092
rect 26424 11086 26476 11092
rect 26160 11070 26280 11086
rect 26252 10810 26280 11070
rect 26332 11008 26384 11014
rect 26332 10950 26384 10956
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26252 10062 26280 10746
rect 26344 10742 26372 10950
rect 26332 10736 26384 10742
rect 26332 10678 26384 10684
rect 26436 10266 26464 11086
rect 27436 11076 27488 11082
rect 27436 11018 27488 11024
rect 27448 10810 27476 11018
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26344 9654 26372 10066
rect 26332 9648 26384 9654
rect 26332 9590 26384 9596
rect 26436 8974 26464 10202
rect 27632 10130 27660 11630
rect 28000 11286 28028 11834
rect 27988 11280 28040 11286
rect 27988 11222 28040 11228
rect 27804 11144 27856 11150
rect 27724 11092 27804 11098
rect 27724 11086 27856 11092
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 27724 11070 27844 11086
rect 27724 10470 27752 11070
rect 27804 11008 27856 11014
rect 27804 10950 27856 10956
rect 27816 10742 27844 10950
rect 27804 10736 27856 10742
rect 27804 10678 27856 10684
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27724 10010 27752 10406
rect 27632 9994 27752 10010
rect 27620 9988 27752 9994
rect 27672 9982 27752 9988
rect 27620 9930 27672 9936
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 26884 9444 26936 9450
rect 26884 9386 26936 9392
rect 26424 8968 26476 8974
rect 26424 8910 26476 8916
rect 26896 8634 26924 9386
rect 27356 9178 27384 9590
rect 27724 9518 27752 9982
rect 27816 9926 27844 10678
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 27908 10266 27936 10610
rect 28092 10606 28120 11086
rect 28080 10600 28132 10606
rect 28080 10542 28132 10548
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 27896 10260 27948 10266
rect 27896 10202 27948 10208
rect 28000 10130 28028 10406
rect 27988 10124 28040 10130
rect 27988 10066 28040 10072
rect 27804 9920 27856 9926
rect 27804 9862 27856 9868
rect 27712 9512 27764 9518
rect 27712 9454 27764 9460
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 26884 8628 26936 8634
rect 26884 8570 26936 8576
rect 28184 8498 28212 12406
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28276 11150 28304 11494
rect 28264 11144 28316 11150
rect 28264 11086 28316 11092
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 26054 7984 26110 7993
rect 26054 7919 26110 7928
rect 28368 7585 28396 29514
rect 28448 16448 28500 16454
rect 28446 16416 28448 16425
rect 28500 16416 28502 16425
rect 28446 16351 28502 16360
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28552 15026 28580 15302
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28644 8906 28672 29514
rect 29460 29504 29512 29510
rect 29460 29446 29512 29452
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29184 29028 29236 29034
rect 29184 28970 29236 28976
rect 29092 28552 29144 28558
rect 29092 28494 29144 28500
rect 29104 28150 29132 28494
rect 29092 28144 29144 28150
rect 29092 28086 29144 28092
rect 28908 27396 28960 27402
rect 28908 27338 28960 27344
rect 28920 27130 28948 27338
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 29104 26994 29132 28086
rect 29092 26988 29144 26994
rect 29092 26930 29144 26936
rect 29000 25900 29052 25906
rect 29000 25842 29052 25848
rect 29012 25498 29040 25842
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 29104 25294 29132 26930
rect 29092 25288 29144 25294
rect 29012 25248 29092 25276
rect 28908 24132 28960 24138
rect 28908 24074 28960 24080
rect 28920 23866 28948 24074
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 29012 23730 29040 25248
rect 29092 25230 29144 25236
rect 29196 23769 29224 28970
rect 29288 28665 29316 29106
rect 29274 28656 29330 28665
rect 29274 28591 29330 28600
rect 29274 27296 29330 27305
rect 29274 27231 29330 27240
rect 29288 27062 29316 27231
rect 29276 27056 29328 27062
rect 29276 26998 29328 27004
rect 29276 26308 29328 26314
rect 29276 26250 29328 26256
rect 29288 25945 29316 26250
rect 29274 25936 29330 25945
rect 29274 25871 29330 25880
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29288 24585 29316 24754
rect 29274 24576 29330 24585
rect 29274 24511 29330 24520
rect 29274 23896 29330 23905
rect 29274 23831 29330 23840
rect 29288 23798 29316 23831
rect 29276 23792 29328 23798
rect 29182 23760 29238 23769
rect 29000 23724 29052 23730
rect 29276 23734 29328 23740
rect 29182 23695 29238 23704
rect 29000 23666 29052 23672
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 28920 22098 28948 22646
rect 29274 22536 29330 22545
rect 29274 22471 29330 22480
rect 28908 22092 28960 22098
rect 28908 22034 28960 22040
rect 29288 22030 29316 22471
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 28816 21616 28868 21622
rect 28816 21558 28868 21564
rect 28828 21146 28856 21558
rect 28816 21140 28868 21146
rect 28816 21082 28868 21088
rect 29012 20942 29040 21966
rect 29184 21888 29236 21894
rect 29184 21830 29236 21836
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 29012 20534 29040 20878
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28920 19514 28948 19722
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 29012 19378 29040 20470
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 29104 18834 29132 20266
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 28908 18352 28960 18358
rect 28908 18294 28960 18300
rect 28920 17882 28948 18294
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28724 17264 28776 17270
rect 28724 17206 28776 17212
rect 28736 16794 28764 17206
rect 28724 16788 28776 16794
rect 28724 16730 28776 16736
rect 29092 16720 29144 16726
rect 29090 16688 29092 16697
rect 29144 16688 29146 16697
rect 29090 16623 29146 16632
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 28920 16182 28948 16390
rect 28908 16176 28960 16182
rect 28908 16118 28960 16124
rect 29092 15496 29144 15502
rect 29092 15438 29144 15444
rect 29104 14482 29132 15438
rect 29092 14476 29144 14482
rect 29092 14418 29144 14424
rect 28908 14340 28960 14346
rect 28908 14282 28960 14288
rect 28920 14074 28948 14282
rect 29196 14278 29224 21830
rect 29274 21176 29330 21185
rect 29274 21111 29330 21120
rect 29288 20942 29316 21111
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 29274 19816 29330 19825
rect 29274 19751 29330 19760
rect 29288 19446 29316 19751
rect 29276 19440 29328 19446
rect 29276 19382 29328 19388
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 29380 18465 29408 18702
rect 29366 18456 29422 18465
rect 29366 18391 29422 18400
rect 29274 17096 29330 17105
rect 29274 17031 29330 17040
rect 29288 16590 29316 17031
rect 29276 16584 29328 16590
rect 29276 16526 29328 16532
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29380 15065 29408 15438
rect 29366 15056 29422 15065
rect 29366 14991 29422 15000
rect 29184 14272 29236 14278
rect 29184 14214 29236 14220
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 28828 12850 28856 13874
rect 29288 13705 29316 13874
rect 29274 13696 29330 13705
rect 29274 13631 29330 13640
rect 28908 13252 28960 13258
rect 28908 13194 28960 13200
rect 28920 12986 28948 13194
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 28816 12844 28868 12850
rect 29276 12844 29328 12850
rect 28868 12804 28948 12832
rect 28816 12786 28868 12792
rect 28920 12238 28948 12804
rect 29276 12786 29328 12792
rect 29288 12345 29316 12786
rect 29274 12336 29330 12345
rect 29274 12271 29330 12280
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 28920 11150 28948 12174
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29012 11354 29040 11698
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 29368 11144 29420 11150
rect 29368 11086 29420 11092
rect 28920 9586 28948 11086
rect 29380 10985 29408 11086
rect 29366 10976 29422 10985
rect 29366 10911 29422 10920
rect 29000 10056 29052 10062
rect 29000 9998 29052 10004
rect 29012 9654 29040 9998
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 29366 9616 29422 9625
rect 28908 9580 28960 9586
rect 29366 9551 29422 9560
rect 28908 9522 28960 9528
rect 29380 9450 29408 9551
rect 29368 9444 29420 9450
rect 29368 9386 29420 9392
rect 28632 8900 28684 8906
rect 28632 8842 28684 8848
rect 29276 8492 29328 8498
rect 29276 8434 29328 8440
rect 29288 8265 29316 8434
rect 29274 8256 29330 8265
rect 29274 8191 29330 8200
rect 29368 7880 29420 7886
rect 29182 7848 29238 7857
rect 29368 7822 29420 7828
rect 29182 7783 29238 7792
rect 29196 7750 29224 7783
rect 29184 7744 29236 7750
rect 29184 7686 29236 7692
rect 29380 7585 29408 7822
rect 28354 7576 28410 7585
rect 28354 7511 28410 7520
rect 29366 7576 29422 7585
rect 29366 7511 29422 7520
rect 29472 7313 29500 29446
rect 29552 26784 29604 26790
rect 29552 26726 29604 26732
rect 29564 7954 29592 26726
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29458 7304 29514 7313
rect 29458 7239 29514 7248
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29104 6322 29132 6598
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29368 6248 29420 6254
rect 29366 6216 29368 6225
rect 29420 6216 29422 6225
rect 29366 6151 29422 6160
rect 29656 5846 29684 19110
rect 29748 7818 29776 30126
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 29736 7812 29788 7818
rect 29736 7754 29788 7760
rect 29840 7342 29868 20742
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29644 5840 29696 5846
rect 29644 5782 29696 5788
rect 29276 5228 29328 5234
rect 29276 5170 29328 5176
rect 29288 4865 29316 5170
rect 29274 4856 29330 4865
rect 29274 4791 29330 4800
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 25332 4282 25360 4558
rect 25320 4276 25372 4282
rect 25320 4218 25372 4224
rect 25044 3936 25096 3942
rect 25044 3878 25096 3884
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 25332 3058 25360 4218
rect 29274 3496 29330 3505
rect 29274 3431 29276 3440
rect 29328 3431 29330 3440
rect 29276 3402 29328 3408
rect 28724 3120 28776 3126
rect 28722 3088 28724 3097
rect 28776 3088 28778 3097
rect 25320 3052 25372 3058
rect 28722 3023 28778 3032
rect 29000 3052 29052 3058
rect 25320 2994 25372 3000
rect 29000 2994 29052 3000
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 24030 2816 24086 2825
rect 24030 2751 24086 2760
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23676 2514 23704 2586
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 24492 2440 24544 2446
rect 25872 2440 25924 2446
rect 24492 2382 24544 2388
rect 25870 2408 25872 2417
rect 25924 2408 25926 2417
rect 23388 2372 23440 2378
rect 23388 2314 23440 2320
rect 24504 800 24532 2382
rect 25780 2372 25832 2378
rect 25870 2343 25926 2352
rect 27068 2372 27120 2378
rect 25780 2314 25832 2320
rect 27068 2314 27120 2320
rect 28356 2372 28408 2378
rect 28356 2314 28408 2320
rect 25792 800 25820 2314
rect 27080 800 27108 2314
rect 27252 2304 27304 2310
rect 27252 2246 27304 2252
rect 28172 2304 28224 2310
rect 28172 2246 28224 2252
rect 27264 1834 27292 2246
rect 28184 2038 28212 2246
rect 28172 2032 28224 2038
rect 28172 1974 28224 1980
rect 27252 1828 27304 1834
rect 27252 1770 27304 1776
rect 28368 800 28396 2314
rect 18 0 74 800
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29012 105 29040 2994
rect 29090 2952 29146 2961
rect 29090 2887 29092 2896
rect 29144 2887 29146 2896
rect 29092 2858 29144 2864
rect 29276 2372 29328 2378
rect 29276 2314 29328 2320
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 29196 1698 29224 2246
rect 29288 2145 29316 2314
rect 29274 2136 29330 2145
rect 29274 2071 29330 2080
rect 29184 1692 29236 1698
rect 29184 1634 29236 1640
rect 29380 785 29408 2994
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 29656 800 29684 2382
rect 29366 776 29422 785
rect 29366 711 29422 720
rect 28998 96 29054 105
rect 28998 31 29054 40
rect 29642 0 29698 800
<< via2 >>
rect 938 32680 994 32736
rect 846 30132 848 30152
rect 848 30132 900 30152
rect 900 30132 902 30152
rect 846 30096 902 30132
rect 29366 32680 29422 32736
rect 1214 31320 1270 31376
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 28538 31320 28594 31376
rect 1398 28600 1454 28656
rect 846 27412 848 27432
rect 848 27412 900 27432
rect 900 27412 902 27432
rect 846 27376 902 27412
rect 1490 25880 1546 25936
rect 846 24656 902 24712
rect 846 23724 902 23760
rect 846 23704 848 23724
rect 848 23704 900 23724
rect 900 23704 902 23724
rect 846 22344 902 22400
rect 1674 21936 1730 21992
rect 846 21256 902 21312
rect 846 19896 902 19952
rect 1674 19796 1676 19816
rect 1676 19796 1728 19816
rect 1728 19796 1730 19816
rect 1674 19760 1730 19796
rect 846 18536 902 18592
rect 846 17212 848 17232
rect 848 17212 900 17232
rect 900 17212 902 17232
rect 846 17176 902 17212
rect 846 16532 848 16552
rect 848 16532 900 16552
rect 900 16532 902 16552
rect 846 16496 902 16532
rect 1490 15000 1546 15056
rect 1398 13640 1454 13696
rect 846 12180 848 12200
rect 848 12180 900 12200
rect 900 12180 902 12200
rect 846 12144 902 12180
rect 846 10784 902 10840
rect 1674 10668 1730 10704
rect 1674 10648 1676 10668
rect 1676 10648 1728 10668
rect 1728 10648 1730 10668
rect 846 7656 902 7712
rect 1398 8200 1454 8256
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 846 4936 902 4992
rect 846 3576 902 3632
rect 2042 7928 2098 7984
rect 2686 22636 2742 22672
rect 2686 22616 2688 22636
rect 2688 22616 2740 22636
rect 2740 22616 2742 22636
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4802 27532 4858 27568
rect 4802 27512 4804 27532
rect 4804 27512 4856 27532
rect 4856 27512 4858 27532
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 5354 23060 5356 23080
rect 5356 23060 5408 23080
rect 5408 23060 5410 23080
rect 5354 23024 5410 23060
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 7102 27396 7158 27432
rect 7102 27376 7104 27396
rect 7104 27376 7156 27396
rect 7156 27376 7158 27396
rect 6182 22616 6238 22672
rect 6366 22636 6422 22672
rect 6366 22616 6368 22636
rect 6368 22616 6420 22636
rect 6420 22616 6422 22636
rect 6090 20884 6092 20904
rect 6092 20884 6144 20904
rect 6144 20884 6146 20904
rect 6090 20848 6146 20884
rect 7746 27512 7802 27568
rect 7654 27276 7656 27296
rect 7656 27276 7708 27296
rect 7708 27276 7710 27296
rect 7654 27240 7710 27276
rect 7838 27396 7894 27432
rect 7838 27376 7840 27396
rect 7840 27376 7892 27396
rect 7892 27376 7894 27396
rect 7470 23060 7472 23080
rect 7472 23060 7524 23080
rect 7524 23060 7526 23080
rect 7470 23024 7526 23060
rect 6550 21836 6552 21856
rect 6552 21836 6604 21856
rect 6604 21836 6606 21856
rect 6550 21800 6606 21836
rect 7746 21800 7802 21856
rect 6826 12824 6882 12880
rect 7930 19660 7932 19680
rect 7932 19660 7984 19680
rect 7984 19660 7986 19680
rect 7930 19624 7986 19660
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1950 5752 2006 5808
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5262 7384 5318 7440
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 6642 9324 6644 9344
rect 6644 9324 6696 9344
rect 6696 9324 6698 9344
rect 6642 9288 6698 9324
rect 7470 9288 7526 9344
rect 7378 7792 7434 7848
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 8482 12844 8538 12880
rect 8482 12824 8484 12844
rect 8484 12824 8536 12844
rect 8536 12824 8538 12844
rect 9586 27240 9642 27296
rect 9770 23724 9826 23760
rect 9770 23704 9772 23724
rect 9772 23704 9824 23724
rect 9824 23704 9826 23724
rect 9770 21664 9826 21720
rect 9218 20304 9274 20360
rect 9402 19372 9458 19408
rect 9402 19352 9404 19372
rect 9404 19352 9456 19372
rect 9456 19352 9458 19372
rect 9126 17856 9182 17912
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4986 2524 4988 2544
rect 4988 2524 5040 2544
rect 5040 2524 5042 2544
rect 4986 2488 5042 2524
rect 938 2080 994 2136
rect 846 856 902 912
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 9678 18844 9680 18864
rect 9680 18844 9732 18864
rect 9732 18844 9734 18864
rect 9678 18808 9734 18844
rect 9678 12180 9680 12200
rect 9680 12180 9732 12200
rect 9732 12180 9734 12200
rect 9678 12144 9734 12180
rect 10322 22344 10378 22400
rect 11150 23740 11152 23760
rect 11152 23740 11204 23760
rect 11204 23740 11206 23760
rect 11150 23704 11206 23740
rect 11426 22344 11482 22400
rect 12530 29008 12586 29064
rect 12254 24148 12256 24168
rect 12256 24148 12308 24168
rect 12308 24148 12310 24168
rect 12254 24112 12310 24148
rect 10230 17448 10286 17504
rect 12070 21664 12126 21720
rect 11702 20576 11758 20632
rect 10046 8336 10102 8392
rect 10322 7928 10378 7984
rect 10690 7284 10692 7304
rect 10692 7284 10744 7304
rect 10744 7284 10746 7304
rect 10690 7248 10746 7284
rect 10322 5652 10324 5672
rect 10324 5652 10376 5672
rect 10376 5652 10378 5672
rect 10322 5616 10378 5652
rect 10414 5208 10470 5264
rect 12622 24112 12678 24168
rect 12254 17448 12310 17504
rect 13174 21664 13230 21720
rect 13818 20576 13874 20632
rect 12806 19352 12862 19408
rect 10966 11756 11022 11792
rect 10966 11736 10968 11756
rect 10968 11736 11020 11756
rect 11020 11736 11022 11756
rect 11150 7928 11206 7984
rect 11150 5908 11206 5944
rect 11150 5888 11152 5908
rect 11152 5888 11204 5908
rect 11204 5888 11206 5908
rect 10966 5652 10968 5672
rect 10968 5652 11020 5672
rect 11020 5652 11022 5672
rect 10966 5616 11022 5652
rect 10966 3476 10968 3496
rect 10968 3476 11020 3496
rect 11020 3476 11022 3496
rect 10966 3440 11022 3476
rect 14370 23724 14426 23760
rect 14370 23704 14372 23724
rect 14372 23704 14424 23724
rect 14424 23704 14426 23724
rect 14186 21972 14188 21992
rect 14188 21972 14240 21992
rect 14240 21972 14242 21992
rect 14186 21936 14242 21972
rect 14462 21800 14518 21856
rect 14186 20304 14242 20360
rect 14922 23704 14978 23760
rect 14646 19252 14648 19272
rect 14648 19252 14700 19272
rect 14700 19252 14702 19272
rect 14646 19216 14702 19252
rect 14002 17856 14058 17912
rect 12622 11736 12678 11792
rect 12714 11636 12716 11656
rect 12716 11636 12768 11656
rect 12768 11636 12770 11656
rect 12714 11600 12770 11636
rect 12898 11328 12954 11384
rect 13082 11328 13138 11384
rect 14094 13776 14150 13832
rect 13818 12144 13874 12200
rect 13910 11600 13966 11656
rect 11610 6296 11666 6352
rect 14094 11600 14150 11656
rect 14830 11600 14886 11656
rect 13726 7928 13782 7984
rect 13266 7248 13322 7304
rect 13082 5652 13084 5672
rect 13084 5652 13136 5672
rect 13136 5652 13138 5672
rect 13082 5616 13138 5652
rect 13542 5228 13598 5264
rect 13542 5208 13544 5228
rect 13544 5208 13596 5228
rect 13596 5208 13598 5228
rect 14002 5888 14058 5944
rect 12162 3440 12218 3496
rect 12070 2644 12126 2680
rect 12070 2624 12072 2644
rect 12072 2624 12124 2644
rect 12124 2624 12126 2644
rect 15014 11736 15070 11792
rect 17406 25236 17408 25256
rect 17408 25236 17460 25256
rect 17460 25236 17462 25256
rect 17406 25200 17462 25236
rect 17038 24520 17094 24576
rect 16946 22480 17002 22536
rect 16854 21392 16910 21448
rect 16118 20304 16174 20360
rect 17682 24556 17684 24576
rect 17684 24556 17736 24576
rect 17736 24556 17738 24576
rect 17682 24520 17738 24556
rect 17038 20340 17040 20360
rect 17040 20340 17092 20360
rect 17092 20340 17094 20360
rect 17038 20304 17094 20340
rect 17038 19488 17094 19544
rect 17498 21392 17554 21448
rect 17682 18808 17738 18864
rect 18050 24520 18106 24576
rect 17866 22516 17868 22536
rect 17868 22516 17920 22536
rect 17920 22516 17922 22536
rect 17866 22480 17922 22516
rect 17866 19488 17922 19544
rect 15290 9560 15346 9616
rect 16762 10668 16818 10704
rect 16762 10648 16764 10668
rect 16764 10648 16816 10668
rect 16816 10648 16818 10668
rect 15014 6316 15070 6352
rect 15014 6296 15016 6316
rect 15016 6296 15068 6316
rect 15068 6296 15070 6316
rect 16762 8336 16818 8392
rect 15750 5652 15752 5672
rect 15752 5652 15804 5672
rect 15804 5652 15806 5672
rect 15750 5616 15806 5652
rect 18970 24520 19026 24576
rect 19706 24520 19762 24576
rect 19154 21956 19210 21992
rect 19154 21936 19156 21956
rect 19156 21936 19208 21956
rect 19208 21936 19210 21956
rect 19246 19896 19302 19952
rect 19522 19760 19578 19816
rect 18326 14476 18382 14512
rect 18326 14456 18328 14476
rect 18328 14456 18380 14476
rect 18380 14456 18382 14476
rect 18602 14476 18658 14512
rect 18602 14456 18604 14476
rect 18604 14456 18656 14476
rect 18656 14456 18658 14476
rect 17222 8336 17278 8392
rect 17590 7520 17646 7576
rect 17774 7248 17830 7304
rect 18510 7248 18566 7304
rect 18878 10668 18934 10704
rect 18878 10648 18880 10668
rect 18880 10648 18932 10668
rect 18932 10648 18934 10668
rect 19614 19624 19670 19680
rect 20074 19896 20130 19952
rect 20166 19760 20222 19816
rect 20074 7404 20130 7440
rect 20074 7384 20076 7404
rect 20076 7384 20128 7404
rect 20128 7384 20130 7404
rect 19982 5752 20038 5808
rect 19338 3596 19394 3632
rect 19338 3576 19340 3596
rect 19340 3576 19392 3596
rect 19392 3576 19394 3596
rect 18878 2252 18880 2272
rect 18880 2252 18932 2272
rect 18932 2252 18934 2272
rect 18878 2216 18934 2252
rect 25226 21936 25282 21992
rect 23478 7384 23534 7440
rect 22006 2760 22062 2816
rect 23110 3576 23166 3632
rect 28906 29960 28962 30016
rect 26054 7928 26110 7984
rect 28446 16396 28448 16416
rect 28448 16396 28500 16416
rect 28500 16396 28502 16416
rect 28446 16360 28502 16396
rect 29274 28600 29330 28656
rect 29274 27240 29330 27296
rect 29274 25880 29330 25936
rect 29274 24520 29330 24576
rect 29274 23840 29330 23896
rect 29182 23704 29238 23760
rect 29274 22480 29330 22536
rect 29090 16668 29092 16688
rect 29092 16668 29144 16688
rect 29144 16668 29146 16688
rect 29090 16632 29146 16668
rect 29274 21120 29330 21176
rect 29274 19760 29330 19816
rect 29366 18400 29422 18456
rect 29274 17040 29330 17096
rect 29366 15000 29422 15056
rect 29274 13640 29330 13696
rect 29274 12280 29330 12336
rect 29366 10920 29422 10976
rect 29366 9560 29422 9616
rect 29274 8200 29330 8256
rect 29182 7792 29238 7848
rect 28354 7520 28410 7576
rect 29366 7520 29422 7576
rect 29458 7248 29514 7304
rect 29366 6196 29368 6216
rect 29368 6196 29420 6216
rect 29420 6196 29422 6216
rect 29366 6160 29422 6196
rect 29274 4800 29330 4856
rect 29274 3460 29330 3496
rect 29274 3440 29276 3460
rect 29276 3440 29328 3460
rect 29328 3440 29330 3460
rect 28722 3068 28724 3088
rect 28724 3068 28776 3088
rect 28776 3068 28778 3088
rect 28722 3032 28778 3068
rect 24030 2760 24086 2816
rect 25870 2388 25872 2408
rect 25872 2388 25924 2408
rect 25924 2388 25926 2408
rect 25870 2352 25926 2388
rect 29090 2916 29146 2952
rect 29090 2896 29092 2916
rect 29092 2896 29144 2916
rect 29144 2896 29146 2916
rect 29274 2080 29330 2136
rect 29366 720 29422 776
rect 28998 40 29054 96
<< metal3 >>
rect 0 32738 800 32768
rect 933 32738 999 32741
rect 0 32736 999 32738
rect 0 32680 938 32736
rect 994 32680 999 32736
rect 0 32678 999 32680
rect 0 32648 800 32678
rect 933 32675 999 32678
rect 29361 32738 29427 32741
rect 30103 32738 30903 32768
rect 29361 32736 30903 32738
rect 29361 32680 29366 32736
rect 29422 32680 30903 32736
rect 29361 32678 30903 32680
rect 29361 32675 29427 32678
rect 30103 32648 30903 32678
rect 0 31378 800 31408
rect 1209 31378 1275 31381
rect 0 31376 1275 31378
rect 0 31320 1214 31376
rect 1270 31320 1275 31376
rect 0 31318 1275 31320
rect 0 31288 800 31318
rect 1209 31315 1275 31318
rect 28533 31378 28599 31381
rect 30103 31378 30903 31408
rect 28533 31376 30903 31378
rect 28533 31320 28538 31376
rect 28594 31320 30903 31376
rect 28533 31318 30903 31320
rect 28533 31315 28599 31318
rect 30103 31288 30903 31318
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 841 30154 907 30157
rect 798 30152 907 30154
rect 798 30096 846 30152
rect 902 30096 907 30152
rect 798 30091 907 30096
rect 798 30048 858 30091
rect 0 29958 858 30048
rect 28901 30018 28967 30021
rect 30103 30018 30903 30048
rect 28901 30016 30903 30018
rect 28901 29960 28906 30016
rect 28962 29960 30903 30016
rect 28901 29958 30903 29960
rect 0 29928 800 29958
rect 28901 29955 28967 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 30103 29928 30903 29958
rect 4210 29887 4526 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 12525 29068 12591 29069
rect 12525 29064 12572 29068
rect 12636 29066 12642 29068
rect 12525 29008 12530 29064
rect 12525 29004 12572 29008
rect 12636 29006 12682 29066
rect 12636 29004 12642 29006
rect 12525 29003 12591 29004
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 0 28658 800 28688
rect 1393 28658 1459 28661
rect 0 28656 1459 28658
rect 0 28600 1398 28656
rect 1454 28600 1459 28656
rect 0 28598 1459 28600
rect 0 28568 800 28598
rect 1393 28595 1459 28598
rect 29269 28658 29335 28661
rect 30103 28658 30903 28688
rect 29269 28656 30903 28658
rect 29269 28600 29274 28656
rect 29330 28600 30903 28656
rect 29269 28598 30903 28600
rect 29269 28595 29335 28598
rect 30103 28568 30903 28598
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 4797 27570 4863 27573
rect 7741 27570 7807 27573
rect 4797 27568 7807 27570
rect 4797 27512 4802 27568
rect 4858 27512 7746 27568
rect 7802 27512 7807 27568
rect 4797 27510 7807 27512
rect 4797 27507 4863 27510
rect 7741 27507 7807 27510
rect 841 27434 907 27437
rect 798 27432 907 27434
rect 798 27376 846 27432
rect 902 27376 907 27432
rect 798 27371 907 27376
rect 7097 27434 7163 27437
rect 7833 27434 7899 27437
rect 7097 27432 7899 27434
rect 7097 27376 7102 27432
rect 7158 27376 7838 27432
rect 7894 27376 7899 27432
rect 7097 27374 7899 27376
rect 7097 27371 7163 27374
rect 7833 27371 7899 27374
rect 798 27328 858 27371
rect 0 27238 858 27328
rect 7649 27298 7715 27301
rect 9581 27298 9647 27301
rect 7649 27296 9647 27298
rect 7649 27240 7654 27296
rect 7710 27240 9586 27296
rect 9642 27240 9647 27296
rect 7649 27238 9647 27240
rect 0 27208 800 27238
rect 7649 27235 7715 27238
rect 9581 27235 9647 27238
rect 29269 27298 29335 27301
rect 30103 27298 30903 27328
rect 29269 27296 30903 27298
rect 29269 27240 29274 27296
rect 29330 27240 30903 27296
rect 29269 27238 30903 27240
rect 29269 27235 29335 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 30103 27208 30903 27238
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 0 25938 800 25968
rect 1485 25938 1551 25941
rect 0 25936 1551 25938
rect 0 25880 1490 25936
rect 1546 25880 1551 25936
rect 0 25878 1551 25880
rect 0 25848 800 25878
rect 1485 25875 1551 25878
rect 29269 25938 29335 25941
rect 30103 25938 30903 25968
rect 29269 25936 30903 25938
rect 29269 25880 29274 25936
rect 29330 25880 30903 25936
rect 29269 25878 30903 25880
rect 29269 25875 29335 25878
rect 30103 25848 30903 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 17401 25258 17467 25261
rect 17718 25258 17724 25260
rect 17401 25256 17724 25258
rect 17401 25200 17406 25256
rect 17462 25200 17724 25256
rect 17401 25198 17724 25200
rect 17401 25195 17467 25198
rect 17718 25196 17724 25198
rect 17788 25196 17794 25260
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 17033 24578 17099 24581
rect 17677 24578 17743 24581
rect 17033 24576 17743 24578
rect 17033 24520 17038 24576
rect 17094 24520 17682 24576
rect 17738 24520 17743 24576
rect 17033 24518 17743 24520
rect 0 24488 800 24518
rect 17033 24515 17099 24518
rect 17677 24515 17743 24518
rect 18045 24578 18111 24581
rect 18965 24578 19031 24581
rect 19701 24578 19767 24581
rect 18045 24576 19767 24578
rect 18045 24520 18050 24576
rect 18106 24520 18970 24576
rect 19026 24520 19706 24576
rect 19762 24520 19767 24576
rect 18045 24518 19767 24520
rect 18045 24515 18111 24518
rect 18965 24515 19031 24518
rect 19701 24515 19767 24518
rect 29269 24578 29335 24581
rect 30103 24578 30903 24608
rect 29269 24576 30903 24578
rect 29269 24520 29274 24576
rect 29330 24520 30903 24576
rect 29269 24518 30903 24520
rect 29269 24515 29335 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 30103 24488 30903 24518
rect 4210 24447 4526 24448
rect 12249 24170 12315 24173
rect 12617 24170 12683 24173
rect 12249 24168 12683 24170
rect 12249 24112 12254 24168
rect 12310 24112 12622 24168
rect 12678 24112 12683 24168
rect 12249 24110 12683 24112
rect 12249 24107 12315 24110
rect 12617 24107 12683 24110
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 29269 23898 29335 23901
rect 30103 23898 30903 23928
rect 0 23808 858 23898
rect 29269 23896 30903 23898
rect 29269 23840 29274 23896
rect 29330 23840 30903 23896
rect 29269 23838 30903 23840
rect 29269 23835 29335 23838
rect 30103 23808 30903 23838
rect 798 23765 858 23808
rect 798 23760 907 23765
rect 798 23704 846 23760
rect 902 23704 907 23760
rect 798 23702 907 23704
rect 841 23699 907 23702
rect 9765 23762 9831 23765
rect 11145 23762 11211 23765
rect 9765 23760 11211 23762
rect 9765 23704 9770 23760
rect 9826 23704 11150 23760
rect 11206 23704 11211 23760
rect 9765 23702 11211 23704
rect 9765 23699 9831 23702
rect 11145 23699 11211 23702
rect 14365 23762 14431 23765
rect 14917 23762 14983 23765
rect 29177 23762 29243 23765
rect 14365 23760 29243 23762
rect 14365 23704 14370 23760
rect 14426 23704 14922 23760
rect 14978 23704 29182 23760
rect 29238 23704 29243 23760
rect 14365 23702 29243 23704
rect 14365 23699 14431 23702
rect 14917 23699 14983 23702
rect 29177 23699 29243 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 5349 23082 5415 23085
rect 7465 23082 7531 23085
rect 5349 23080 7531 23082
rect 5349 23024 5354 23080
rect 5410 23024 7470 23080
rect 7526 23024 7531 23080
rect 5349 23022 7531 23024
rect 5349 23019 5415 23022
rect 7465 23019 7531 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 2681 22674 2747 22677
rect 6177 22674 6243 22677
rect 6361 22674 6427 22677
rect 2681 22672 6427 22674
rect 2681 22616 2686 22672
rect 2742 22616 6182 22672
rect 6238 22616 6366 22672
rect 6422 22616 6427 22672
rect 2681 22614 6427 22616
rect 2681 22611 2747 22614
rect 6177 22611 6243 22614
rect 6361 22611 6427 22614
rect 0 22538 800 22568
rect 16941 22538 17007 22541
rect 17861 22538 17927 22541
rect 0 22448 858 22538
rect 16941 22536 17927 22538
rect 16941 22480 16946 22536
rect 17002 22480 17866 22536
rect 17922 22480 17927 22536
rect 16941 22478 17927 22480
rect 16941 22475 17007 22478
rect 17861 22475 17927 22478
rect 29269 22538 29335 22541
rect 30103 22538 30903 22568
rect 29269 22536 30903 22538
rect 29269 22480 29274 22536
rect 29330 22480 30903 22536
rect 29269 22478 30903 22480
rect 29269 22475 29335 22478
rect 30103 22448 30903 22478
rect 798 22405 858 22448
rect 798 22400 907 22405
rect 798 22344 846 22400
rect 902 22344 907 22400
rect 798 22342 907 22344
rect 841 22339 907 22342
rect 10317 22402 10383 22405
rect 11421 22402 11487 22405
rect 10317 22400 11487 22402
rect 10317 22344 10322 22400
rect 10378 22344 11426 22400
rect 11482 22344 11487 22400
rect 10317 22342 11487 22344
rect 10317 22339 10383 22342
rect 11421 22339 11487 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 1669 21994 1735 21997
rect 1669 21992 12450 21994
rect 1669 21936 1674 21992
rect 1730 21936 12450 21992
rect 1669 21934 12450 21936
rect 1669 21931 1735 21934
rect 6545 21858 6611 21861
rect 7741 21858 7807 21861
rect 6545 21856 7807 21858
rect 6545 21800 6550 21856
rect 6606 21800 7746 21856
rect 7802 21800 7807 21856
rect 6545 21798 7807 21800
rect 12390 21858 12450 21934
rect 12566 21932 12572 21996
rect 12636 21994 12642 21996
rect 14181 21994 14247 21997
rect 12636 21992 14247 21994
rect 12636 21936 14186 21992
rect 14242 21936 14247 21992
rect 12636 21934 14247 21936
rect 12636 21932 12642 21934
rect 14181 21931 14247 21934
rect 19149 21994 19215 21997
rect 25221 21994 25287 21997
rect 19149 21992 25287 21994
rect 19149 21936 19154 21992
rect 19210 21936 25226 21992
rect 25282 21936 25287 21992
rect 19149 21934 25287 21936
rect 19149 21931 19215 21934
rect 25221 21931 25287 21934
rect 14457 21858 14523 21861
rect 12390 21856 14523 21858
rect 12390 21800 14462 21856
rect 14518 21800 14523 21856
rect 12390 21798 14523 21800
rect 6545 21795 6611 21798
rect 7741 21795 7807 21798
rect 14457 21795 14523 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 9765 21722 9831 21725
rect 12065 21722 12131 21725
rect 13169 21722 13235 21725
rect 9765 21720 13235 21722
rect 9765 21664 9770 21720
rect 9826 21664 12070 21720
rect 12126 21664 13174 21720
rect 13230 21664 13235 21720
rect 9765 21662 13235 21664
rect 9765 21659 9831 21662
rect 12065 21659 12131 21662
rect 13169 21659 13235 21662
rect 16849 21450 16915 21453
rect 16982 21450 16988 21452
rect 16849 21448 16988 21450
rect 16849 21392 16854 21448
rect 16910 21392 16988 21448
rect 16849 21390 16988 21392
rect 16849 21387 16915 21390
rect 16982 21388 16988 21390
rect 17052 21450 17058 21452
rect 17493 21450 17559 21453
rect 17052 21448 17559 21450
rect 17052 21392 17498 21448
rect 17554 21392 17559 21448
rect 17052 21390 17559 21392
rect 17052 21388 17058 21390
rect 17493 21387 17559 21390
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 29269 21178 29335 21181
rect 30103 21178 30903 21208
rect 29269 21176 30903 21178
rect 29269 21120 29274 21176
rect 29330 21120 30903 21176
rect 29269 21118 30903 21120
rect 0 21088 800 21118
rect 29269 21115 29335 21118
rect 30103 21088 30903 21118
rect 6085 20908 6151 20909
rect 6085 20906 6132 20908
rect 6040 20904 6132 20906
rect 6040 20848 6090 20904
rect 6040 20846 6132 20848
rect 6085 20844 6132 20846
rect 6196 20844 6202 20908
rect 6085 20843 6151 20844
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 11697 20634 11763 20637
rect 13813 20634 13879 20637
rect 11697 20632 13879 20634
rect 11697 20576 11702 20632
rect 11758 20576 13818 20632
rect 13874 20576 13879 20632
rect 11697 20574 13879 20576
rect 11697 20571 11763 20574
rect 13813 20571 13879 20574
rect 9213 20364 9279 20365
rect 14181 20364 14247 20365
rect 9213 20362 9260 20364
rect 9168 20360 9260 20362
rect 9168 20304 9218 20360
rect 9168 20302 9260 20304
rect 9213 20300 9260 20302
rect 9324 20300 9330 20364
rect 14181 20362 14228 20364
rect 14136 20360 14228 20362
rect 14292 20362 14298 20364
rect 16113 20362 16179 20365
rect 17033 20362 17099 20365
rect 14292 20360 17099 20362
rect 14136 20304 14186 20360
rect 14292 20304 16118 20360
rect 16174 20304 17038 20360
rect 17094 20304 17099 20360
rect 14136 20302 14228 20304
rect 14181 20300 14228 20302
rect 14292 20302 17099 20304
rect 14292 20300 14298 20302
rect 9213 20299 9279 20300
rect 14181 20299 14247 20300
rect 16113 20299 16179 20302
rect 17033 20299 17099 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 19241 19954 19307 19957
rect 20069 19954 20135 19957
rect 19241 19952 20135 19954
rect 19241 19896 19246 19952
rect 19302 19896 20074 19952
rect 20130 19896 20135 19952
rect 19241 19894 20135 19896
rect 19241 19891 19307 19894
rect 20069 19891 20135 19894
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 1669 19818 1735 19821
rect 19517 19818 19583 19821
rect 20161 19818 20227 19821
rect 1669 19816 20227 19818
rect 1669 19760 1674 19816
rect 1730 19760 19522 19816
rect 19578 19760 20166 19816
rect 20222 19760 20227 19816
rect 1669 19758 20227 19760
rect 0 19728 800 19758
rect 1669 19755 1735 19758
rect 19517 19755 19583 19758
rect 20161 19755 20227 19758
rect 29269 19818 29335 19821
rect 30103 19818 30903 19848
rect 29269 19816 30903 19818
rect 29269 19760 29274 19816
rect 29330 19760 30903 19816
rect 29269 19758 30903 19760
rect 29269 19755 29335 19758
rect 30103 19728 30903 19758
rect 7925 19682 7991 19685
rect 19609 19682 19675 19685
rect 7925 19680 19675 19682
rect 7925 19624 7930 19680
rect 7986 19624 19614 19680
rect 19670 19624 19675 19680
rect 7925 19622 19675 19624
rect 7925 19619 7991 19622
rect 19609 19619 19675 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 17033 19546 17099 19549
rect 17861 19546 17927 19549
rect 17033 19544 17927 19546
rect 17033 19488 17038 19544
rect 17094 19488 17866 19544
rect 17922 19488 17927 19544
rect 17033 19486 17927 19488
rect 17033 19483 17099 19486
rect 17861 19483 17927 19486
rect 9397 19410 9463 19413
rect 12801 19410 12867 19413
rect 9397 19408 12867 19410
rect 9397 19352 9402 19408
rect 9458 19352 12806 19408
rect 12862 19352 12867 19408
rect 9397 19350 12867 19352
rect 9397 19347 9463 19350
rect 12801 19347 12867 19350
rect 14641 19274 14707 19277
rect 14774 19274 14780 19276
rect 14641 19272 14780 19274
rect 14641 19216 14646 19272
rect 14702 19216 14780 19272
rect 14641 19214 14780 19216
rect 14641 19211 14707 19214
rect 14774 19212 14780 19214
rect 14844 19212 14850 19276
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 9673 18866 9739 18869
rect 17677 18868 17743 18869
rect 9806 18866 9812 18868
rect 9673 18864 9812 18866
rect 9673 18808 9678 18864
rect 9734 18808 9812 18864
rect 9673 18806 9812 18808
rect 9673 18803 9739 18806
rect 9806 18804 9812 18806
rect 9876 18804 9882 18868
rect 17677 18864 17724 18868
rect 17788 18866 17794 18868
rect 17677 18808 17682 18864
rect 17677 18804 17724 18808
rect 17788 18806 17834 18866
rect 17788 18804 17794 18806
rect 17677 18803 17743 18804
rect 841 18594 907 18597
rect 798 18592 907 18594
rect 798 18536 846 18592
rect 902 18536 907 18592
rect 798 18531 907 18536
rect 798 18488 858 18531
rect 0 18398 858 18488
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 29361 18458 29427 18461
rect 30103 18458 30903 18488
rect 29361 18456 30903 18458
rect 29361 18400 29366 18456
rect 29422 18400 30903 18456
rect 29361 18398 30903 18400
rect 0 18368 800 18398
rect 29361 18395 29427 18398
rect 30103 18368 30903 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 9121 17914 9187 17917
rect 13997 17914 14063 17917
rect 9121 17912 14063 17914
rect 9121 17856 9126 17912
rect 9182 17856 14002 17912
rect 14058 17856 14063 17912
rect 9121 17854 14063 17856
rect 9121 17851 9187 17854
rect 10225 17506 10291 17509
rect 12249 17506 12315 17509
rect 10225 17504 12315 17506
rect 10225 17448 10230 17504
rect 10286 17448 12254 17504
rect 12310 17448 12315 17504
rect 10225 17446 12315 17448
rect 10225 17443 10291 17446
rect 12249 17443 12315 17446
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 841 17234 907 17237
rect 798 17232 907 17234
rect 798 17176 846 17232
rect 902 17176 907 17232
rect 798 17171 907 17176
rect 798 17128 858 17171
rect 0 17038 858 17128
rect 0 17008 800 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 12390 16690 12450 17854
rect 13997 17851 14063 17854
rect 29269 17098 29335 17101
rect 30103 17098 30903 17128
rect 29269 17096 30903 17098
rect 29269 17040 29274 17096
rect 29330 17040 30903 17096
rect 29269 17038 30903 17040
rect 29269 17035 29335 17038
rect 30103 17008 30903 17038
rect 29085 16690 29151 16693
rect 12390 16688 29151 16690
rect 12390 16632 29090 16688
rect 29146 16632 29151 16688
rect 12390 16630 29151 16632
rect 29085 16627 29151 16630
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 28441 16418 28507 16421
rect 30103 16418 30903 16448
rect 28441 16416 30903 16418
rect 28441 16360 28446 16416
rect 28502 16360 30903 16416
rect 28441 16358 30903 16360
rect 0 16328 800 16358
rect 28441 16355 28507 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 30103 16328 30903 16358
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 29361 15058 29427 15061
rect 30103 15058 30903 15088
rect 29361 15056 30903 15058
rect 29361 15000 29366 15056
rect 29422 15000 30903 15056
rect 29361 14998 30903 15000
rect 29361 14995 29427 14998
rect 30103 14968 30903 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 18321 14514 18387 14517
rect 18597 14514 18663 14517
rect 18321 14512 18663 14514
rect 18321 14456 18326 14512
rect 18382 14456 18602 14512
rect 18658 14456 18663 14512
rect 18321 14454 18663 14456
rect 18321 14451 18387 14454
rect 18597 14451 18663 14454
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 14089 13834 14155 13837
rect 14406 13834 14412 13836
rect 14089 13832 14412 13834
rect 14089 13776 14094 13832
rect 14150 13776 14412 13832
rect 14089 13774 14412 13776
rect 14089 13771 14155 13774
rect 14406 13772 14412 13774
rect 14476 13772 14482 13836
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 29269 13698 29335 13701
rect 30103 13698 30903 13728
rect 29269 13696 30903 13698
rect 29269 13640 29274 13696
rect 29330 13640 30903 13696
rect 29269 13638 30903 13640
rect 29269 13635 29335 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 30103 13608 30903 13638
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 6821 12882 6887 12885
rect 8477 12882 8543 12885
rect 6821 12880 8543 12882
rect 6821 12824 6826 12880
rect 6882 12824 8482 12880
rect 8538 12824 8543 12880
rect 6821 12822 8543 12824
rect 6821 12819 6887 12822
rect 8477 12819 8543 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 29269 12338 29335 12341
rect 30103 12338 30903 12368
rect 0 12248 858 12338
rect 29269 12336 30903 12338
rect 29269 12280 29274 12336
rect 29330 12280 30903 12336
rect 29269 12278 30903 12280
rect 29269 12275 29335 12278
rect 30103 12248 30903 12278
rect 798 12205 858 12248
rect 798 12200 907 12205
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12142 907 12144
rect 841 12139 907 12142
rect 9673 12202 9739 12205
rect 13813 12202 13879 12205
rect 9673 12200 13879 12202
rect 9673 12144 9678 12200
rect 9734 12144 13818 12200
rect 13874 12144 13879 12200
rect 9673 12142 13879 12144
rect 9673 12139 9739 12142
rect 13813 12139 13879 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 10961 11794 11027 11797
rect 12617 11794 12683 11797
rect 15009 11794 15075 11797
rect 10961 11792 15075 11794
rect 10961 11736 10966 11792
rect 11022 11736 12622 11792
rect 12678 11736 15014 11792
rect 15070 11736 15075 11792
rect 10961 11734 15075 11736
rect 10961 11731 11027 11734
rect 12617 11731 12683 11734
rect 15009 11731 15075 11734
rect 12709 11658 12775 11661
rect 13905 11658 13971 11661
rect 14089 11658 14155 11661
rect 14825 11658 14891 11661
rect 12709 11656 14891 11658
rect 12709 11600 12714 11656
rect 12770 11600 13910 11656
rect 13966 11600 14094 11656
rect 14150 11600 14830 11656
rect 14886 11600 14891 11656
rect 12709 11598 14891 11600
rect 12709 11595 12775 11598
rect 13905 11595 13971 11598
rect 14089 11595 14155 11598
rect 14825 11595 14891 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12893 11386 12959 11389
rect 13077 11386 13143 11389
rect 12893 11384 13143 11386
rect 12893 11328 12898 11384
rect 12954 11328 13082 11384
rect 13138 11328 13143 11384
rect 12893 11326 13143 11328
rect 12893 11323 12959 11326
rect 13077 11323 13143 11326
rect 0 10978 800 11008
rect 29361 10978 29427 10981
rect 30103 10978 30903 11008
rect 0 10888 858 10978
rect 29361 10976 30903 10978
rect 29361 10920 29366 10976
rect 29422 10920 30903 10976
rect 29361 10918 30903 10920
rect 29361 10915 29427 10918
rect 798 10845 858 10888
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 30103 10888 30903 10918
rect 4870 10847 5186 10848
rect 798 10840 907 10845
rect 798 10784 846 10840
rect 902 10784 907 10840
rect 798 10782 907 10784
rect 841 10779 907 10782
rect 1669 10706 1735 10709
rect 6126 10706 6132 10708
rect 1669 10704 6132 10706
rect 1669 10648 1674 10704
rect 1730 10648 6132 10704
rect 1669 10646 6132 10648
rect 1669 10643 1735 10646
rect 6126 10644 6132 10646
rect 6196 10644 6202 10708
rect 16757 10706 16823 10709
rect 18873 10706 18939 10709
rect 16757 10704 18939 10706
rect 16757 10648 16762 10704
rect 16818 10648 18878 10704
rect 18934 10648 18939 10704
rect 16757 10646 18939 10648
rect 16757 10643 16823 10646
rect 18873 10643 18939 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 15285 9618 15351 9621
rect 0 9616 15351 9618
rect 0 9560 15290 9616
rect 15346 9560 15351 9616
rect 0 9558 15351 9560
rect 0 9528 800 9558
rect 15285 9555 15351 9558
rect 29361 9618 29427 9621
rect 30103 9618 30903 9648
rect 29361 9616 30903 9618
rect 29361 9560 29366 9616
rect 29422 9560 30903 9616
rect 29361 9558 30903 9560
rect 29361 9555 29427 9558
rect 30103 9528 30903 9558
rect 6637 9346 6703 9349
rect 7465 9346 7531 9349
rect 6637 9344 7531 9346
rect 6637 9288 6642 9344
rect 6698 9288 7470 9344
rect 7526 9288 7531 9344
rect 6637 9286 7531 9288
rect 6637 9283 6703 9286
rect 7465 9283 7531 9286
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 10041 8394 10107 8397
rect 16757 8394 16823 8397
rect 17217 8394 17283 8397
rect 10041 8392 17283 8394
rect 10041 8336 10046 8392
rect 10102 8336 16762 8392
rect 16818 8336 17222 8392
rect 17278 8336 17283 8392
rect 10041 8334 17283 8336
rect 10041 8331 10107 8334
rect 16757 8331 16823 8334
rect 17217 8331 17283 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 29269 8258 29335 8261
rect 30103 8258 30903 8288
rect 29269 8256 30903 8258
rect 29269 8200 29274 8256
rect 29330 8200 30903 8256
rect 29269 8198 30903 8200
rect 29269 8195 29335 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 30103 8168 30903 8198
rect 4210 8127 4526 8128
rect 2037 7986 2103 7989
rect 10317 7986 10383 7989
rect 2037 7984 10383 7986
rect 2037 7928 2042 7984
rect 2098 7928 10322 7984
rect 10378 7928 10383 7984
rect 2037 7926 10383 7928
rect 2037 7923 2103 7926
rect 10317 7923 10383 7926
rect 11145 7986 11211 7989
rect 13721 7986 13787 7989
rect 26049 7986 26115 7989
rect 11145 7984 26115 7986
rect 11145 7928 11150 7984
rect 11206 7928 13726 7984
rect 13782 7928 26054 7984
rect 26110 7928 26115 7984
rect 11145 7926 26115 7928
rect 11145 7923 11211 7926
rect 13721 7923 13787 7926
rect 26049 7923 26115 7926
rect 7373 7850 7439 7853
rect 29177 7850 29243 7853
rect 7373 7848 29243 7850
rect 7373 7792 7378 7848
rect 7434 7792 29182 7848
rect 29238 7792 29243 7848
rect 7373 7790 29243 7792
rect 7373 7787 7439 7790
rect 29177 7787 29243 7790
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 17585 7578 17651 7581
rect 28349 7578 28415 7581
rect 17585 7576 28415 7578
rect 17585 7520 17590 7576
rect 17646 7520 28354 7576
rect 28410 7520 28415 7576
rect 17585 7518 28415 7520
rect 0 7488 800 7518
rect 17585 7515 17651 7518
rect 28349 7515 28415 7518
rect 29361 7578 29427 7581
rect 30103 7578 30903 7608
rect 29361 7576 30903 7578
rect 29361 7520 29366 7576
rect 29422 7520 30903 7576
rect 29361 7518 30903 7520
rect 29361 7515 29427 7518
rect 30103 7488 30903 7518
rect 5257 7442 5323 7445
rect 20069 7442 20135 7445
rect 23473 7442 23539 7445
rect 5257 7440 23539 7442
rect 5257 7384 5262 7440
rect 5318 7384 20074 7440
rect 20130 7384 23478 7440
rect 23534 7384 23539 7440
rect 5257 7382 23539 7384
rect 5257 7379 5323 7382
rect 20069 7379 20135 7382
rect 23473 7379 23539 7382
rect 10685 7306 10751 7309
rect 13261 7306 13327 7309
rect 10685 7304 13327 7306
rect 10685 7248 10690 7304
rect 10746 7248 13266 7304
rect 13322 7248 13327 7304
rect 10685 7246 13327 7248
rect 10685 7243 10751 7246
rect 13261 7243 13327 7246
rect 17769 7306 17835 7309
rect 18505 7306 18571 7309
rect 29453 7306 29519 7309
rect 17769 7304 29519 7306
rect 17769 7248 17774 7304
rect 17830 7248 18510 7304
rect 18566 7248 29458 7304
rect 29514 7248 29519 7304
rect 17769 7246 29519 7248
rect 17769 7243 17835 7246
rect 18505 7243 18571 7246
rect 29453 7243 29519 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 11605 6354 11671 6357
rect 15009 6354 15075 6357
rect 11605 6352 15075 6354
rect 11605 6296 11610 6352
rect 11666 6296 15014 6352
rect 15070 6296 15075 6352
rect 11605 6294 15075 6296
rect 11605 6291 11671 6294
rect 15009 6291 15075 6294
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 29361 6218 29427 6221
rect 30103 6218 30903 6248
rect 29361 6216 30903 6218
rect 29361 6160 29366 6216
rect 29422 6160 30903 6216
rect 29361 6158 30903 6160
rect 0 6128 800 6158
rect 29361 6155 29427 6158
rect 30103 6128 30903 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 11145 5946 11211 5949
rect 13997 5946 14063 5949
rect 11145 5944 14063 5946
rect 11145 5888 11150 5944
rect 11206 5888 14002 5944
rect 14058 5888 14063 5944
rect 11145 5886 14063 5888
rect 11145 5883 11211 5886
rect 13997 5883 14063 5886
rect 1945 5810 2011 5813
rect 19977 5810 20043 5813
rect 1945 5808 20043 5810
rect 1945 5752 1950 5808
rect 2006 5752 19982 5808
rect 20038 5752 20043 5808
rect 1945 5750 20043 5752
rect 1945 5747 2011 5750
rect 19977 5747 20043 5750
rect 10317 5674 10383 5677
rect 10961 5674 11027 5677
rect 10317 5672 11027 5674
rect 10317 5616 10322 5672
rect 10378 5616 10966 5672
rect 11022 5616 11027 5672
rect 10317 5614 11027 5616
rect 10317 5611 10383 5614
rect 10961 5611 11027 5614
rect 13077 5674 13143 5677
rect 15745 5674 15811 5677
rect 13077 5672 15811 5674
rect 13077 5616 13082 5672
rect 13138 5616 15750 5672
rect 15806 5616 15811 5672
rect 13077 5614 15811 5616
rect 13077 5611 13143 5614
rect 15745 5611 15811 5614
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 10409 5266 10475 5269
rect 13537 5266 13603 5269
rect 10409 5264 13603 5266
rect 10409 5208 10414 5264
rect 10470 5208 13542 5264
rect 13598 5208 13603 5264
rect 10409 5206 13603 5208
rect 10409 5203 10475 5206
rect 13537 5203 13603 5206
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 29269 4858 29335 4861
rect 30103 4858 30903 4888
rect 29269 4856 30903 4858
rect 29269 4800 29274 4856
rect 29330 4800 30903 4856
rect 29269 4798 30903 4800
rect 0 4768 800 4798
rect 29269 4795 29335 4798
rect 30103 4768 30903 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 841 3634 907 3637
rect 798 3632 907 3634
rect 798 3576 846 3632
rect 902 3576 907 3632
rect 798 3571 907 3576
rect 19333 3634 19399 3637
rect 23105 3634 23171 3637
rect 19333 3632 23171 3634
rect 19333 3576 19338 3632
rect 19394 3576 23110 3632
rect 23166 3576 23171 3632
rect 19333 3574 23171 3576
rect 19333 3571 19399 3574
rect 23105 3571 23171 3574
rect 798 3528 858 3571
rect 0 3438 858 3528
rect 10961 3498 11027 3501
rect 12157 3498 12223 3501
rect 10961 3496 12223 3498
rect 10961 3440 10966 3496
rect 11022 3440 12162 3496
rect 12218 3440 12223 3496
rect 10961 3438 12223 3440
rect 0 3408 800 3438
rect 10961 3435 11027 3438
rect 12157 3435 12223 3438
rect 29269 3498 29335 3501
rect 30103 3498 30903 3528
rect 29269 3496 30903 3498
rect 29269 3440 29274 3496
rect 29330 3440 30903 3496
rect 29269 3438 30903 3440
rect 29269 3435 29335 3438
rect 30103 3408 30903 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 16982 3028 16988 3092
rect 17052 3090 17058 3092
rect 28717 3090 28783 3093
rect 17052 3088 28783 3090
rect 17052 3032 28722 3088
rect 28778 3032 28783 3088
rect 17052 3030 28783 3032
rect 17052 3028 17058 3030
rect 28717 3027 28783 3030
rect 9254 2892 9260 2956
rect 9324 2954 9330 2956
rect 29085 2954 29151 2957
rect 9324 2952 29151 2954
rect 9324 2896 29090 2952
rect 29146 2896 29151 2952
rect 9324 2894 29151 2896
rect 9324 2892 9330 2894
rect 29085 2891 29151 2894
rect 22001 2818 22067 2821
rect 24025 2818 24091 2821
rect 22001 2816 24091 2818
rect 22001 2760 22006 2816
rect 22062 2760 24030 2816
rect 24086 2760 24091 2816
rect 22001 2758 24091 2760
rect 22001 2755 22067 2758
rect 24025 2755 24091 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12065 2682 12131 2685
rect 14222 2682 14228 2684
rect 12065 2680 14228 2682
rect 12065 2624 12070 2680
rect 12126 2624 14228 2680
rect 12065 2622 14228 2624
rect 12065 2619 12131 2622
rect 14222 2620 14228 2622
rect 14292 2620 14298 2684
rect 4981 2546 5047 2549
rect 14774 2546 14780 2548
rect 4981 2544 14780 2546
rect 4981 2488 4986 2544
rect 5042 2488 14780 2544
rect 4981 2486 14780 2488
rect 4981 2483 5047 2486
rect 14774 2484 14780 2486
rect 14844 2484 14850 2548
rect 14406 2348 14412 2412
rect 14476 2410 14482 2412
rect 25865 2410 25931 2413
rect 14476 2408 25931 2410
rect 14476 2352 25870 2408
rect 25926 2352 25931 2408
rect 14476 2350 25931 2352
rect 14476 2348 14482 2350
rect 25865 2347 25931 2350
rect 9806 2212 9812 2276
rect 9876 2274 9882 2276
rect 18873 2274 18939 2277
rect 9876 2272 18939 2274
rect 9876 2216 18878 2272
rect 18934 2216 18939 2272
rect 9876 2214 18939 2216
rect 9876 2212 9882 2214
rect 18873 2211 18939 2214
rect 4870 2208 5186 2209
rect 0 2138 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 933 2138 999 2141
rect 0 2136 999 2138
rect 0 2080 938 2136
rect 994 2080 999 2136
rect 0 2078 999 2080
rect 0 2048 800 2078
rect 933 2075 999 2078
rect 29269 2138 29335 2141
rect 30103 2138 30903 2168
rect 29269 2136 30903 2138
rect 29269 2080 29274 2136
rect 29330 2080 30903 2136
rect 29269 2078 30903 2080
rect 29269 2075 29335 2078
rect 30103 2048 30903 2078
rect 841 914 907 917
rect 798 912 907 914
rect 798 856 846 912
rect 902 856 907 912
rect 798 851 907 856
rect 798 808 858 851
rect 0 718 858 808
rect 29361 778 29427 781
rect 30103 778 30903 808
rect 29361 776 30903 778
rect 29361 720 29366 776
rect 29422 720 30903 776
rect 29361 718 30903 720
rect 0 688 800 718
rect 29361 715 29427 718
rect 30103 688 30903 718
rect 28993 98 29059 101
rect 30103 98 30903 128
rect 28993 96 30903 98
rect 28993 40 28998 96
rect 29054 40 30903 96
rect 28993 38 30903 40
rect 28993 35 29059 38
rect 30103 8 30903 38
<< via3 >>
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 12572 29064 12636 29068
rect 12572 29008 12586 29064
rect 12586 29008 12636 29064
rect 12572 29004 12636 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 17724 25196 17788 25260
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 12572 21932 12636 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 16988 21388 17052 21452
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 6132 20904 6196 20908
rect 6132 20848 6146 20904
rect 6146 20848 6196 20904
rect 6132 20844 6196 20848
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 9260 20360 9324 20364
rect 9260 20304 9274 20360
rect 9274 20304 9324 20360
rect 9260 20300 9324 20304
rect 14228 20360 14292 20364
rect 14228 20304 14242 20360
rect 14242 20304 14292 20360
rect 14228 20300 14292 20304
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 14780 19212 14844 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 9812 18804 9876 18868
rect 17724 18864 17788 18868
rect 17724 18808 17738 18864
rect 17738 18808 17788 18864
rect 17724 18804 17788 18808
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 14412 13772 14476 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 6132 10644 6196 10708
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 16988 3028 17052 3092
rect 9260 2892 9324 2956
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 14228 2620 14292 2684
rect 14780 2484 14844 2548
rect 14412 2348 14476 2412
rect 9812 2212 9876 2276
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 29952 4528 30512
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 30496 5188 30512
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 12571 29068 12637 29069
rect 12571 29004 12572 29068
rect 12636 29004 12637 29068
rect 12571 29003 12637 29004
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 12574 21997 12634 29003
rect 17723 25260 17789 25261
rect 17723 25196 17724 25260
rect 17788 25196 17789 25260
rect 17723 25195 17789 25196
rect 12571 21996 12637 21997
rect 12571 21932 12572 21996
rect 12636 21932 12637 21996
rect 12571 21931 12637 21932
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 16987 21452 17053 21453
rect 16987 21388 16988 21452
rect 17052 21388 17053 21452
rect 16987 21387 17053 21388
rect 6131 20908 6197 20909
rect 6131 20844 6132 20908
rect 6196 20844 6197 20908
rect 6131 20843 6197 20844
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 6134 10709 6194 20843
rect 9259 20364 9325 20365
rect 9259 20300 9260 20364
rect 9324 20300 9325 20364
rect 9259 20299 9325 20300
rect 14227 20364 14293 20365
rect 14227 20300 14228 20364
rect 14292 20300 14293 20364
rect 14227 20299 14293 20300
rect 6131 10708 6197 10709
rect 6131 10644 6132 10708
rect 6196 10644 6197 10708
rect 6131 10643 6197 10644
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 9262 2957 9322 20299
rect 9811 18868 9877 18869
rect 9811 18804 9812 18868
rect 9876 18804 9877 18868
rect 9811 18803 9877 18804
rect 9259 2956 9325 2957
rect 9259 2892 9260 2956
rect 9324 2892 9325 2956
rect 9259 2891 9325 2892
rect 9814 2277 9874 18803
rect 14230 2685 14290 20299
rect 14779 19276 14845 19277
rect 14779 19212 14780 19276
rect 14844 19212 14845 19276
rect 14779 19211 14845 19212
rect 14411 13836 14477 13837
rect 14411 13772 14412 13836
rect 14476 13772 14477 13836
rect 14411 13771 14477 13772
rect 14227 2684 14293 2685
rect 14227 2620 14228 2684
rect 14292 2620 14293 2684
rect 14227 2619 14293 2620
rect 14414 2413 14474 13771
rect 14782 2549 14842 19211
rect 16990 3093 17050 21387
rect 17726 18869 17786 25195
rect 17723 18868 17789 18869
rect 17723 18804 17724 18868
rect 17788 18804 17789 18868
rect 17723 18803 17789 18804
rect 16987 3092 17053 3093
rect 16987 3028 16988 3092
rect 17052 3028 17053 3092
rect 16987 3027 17053 3028
rect 14779 2548 14845 2549
rect 14779 2484 14780 2548
rect 14844 2484 14845 2548
rect 14779 2483 14845 2484
rect 14411 2412 14477 2413
rect 14411 2348 14412 2412
rect 14476 2348 14477 2412
rect 14411 2347 14477 2348
rect 9811 2276 9877 2277
rect 9811 2212 9812 2276
rect 9876 2212 9877 2276
rect 9811 2211 9877 2212
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0942_
timestamp -3599
transform -1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp -3599
transform -1 0 21436 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp -3599
transform -1 0 22908 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp -3599
transform -1 0 21160 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp -3599
transform -1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp -3599
transform 1 0 18492 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp -3599
transform -1 0 15640 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0949_
timestamp -3599
transform -1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0950_
timestamp -3599
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp -3599
transform -1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp -3599
transform 1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp -3599
transform 1 0 7268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp -3599
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp -3599
transform -1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0956_
timestamp -3599
transform 1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp -3599
transform 1 0 8280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp -3599
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp -3599
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp -3599
transform 1 0 8740 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp -3599
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0962_
timestamp -3599
transform 1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp -3599
transform 1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp -3599
transform -1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0965_
timestamp -3599
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp -3599
transform -1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp -3599
transform 1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp -3599
transform 1 0 19964 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp -3599
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp -3599
transform 1 0 22632 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp -3599
transform 1 0 24472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp -3599
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp -3599
transform -1 0 26128 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0974_
timestamp -3599
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp -3599
transform -1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp -3599
transform 1 0 18492 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp -3599
transform -1 0 18400 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp -3599
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp -3599
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp -3599
transform 1 0 14628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0981_
timestamp -3599
transform 1 0 12788 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp -3599
transform -1 0 13616 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp -3599
transform 1 0 11592 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp -3599
transform -1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp -3599
transform -1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp -3599
transform -1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0987_
timestamp -3599
transform -1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp -3599
transform 1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp -3599
transform 1 0 16192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp -3599
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp -3599
transform -1 0 25760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp -3599
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0993_
timestamp -3599
transform -1 0 19320 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp -3599
transform -1 0 19964 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp -3599
transform 1 0 19780 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp -3599
transform 1 0 17572 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp -3599
transform -1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp -3599
transform -1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0999_
timestamp -3599
transform -1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp -3599
transform 1 0 14076 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp -3599
transform 1 0 13248 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp -3599
transform -1 0 10120 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp -3599
transform -1 0 8740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp -3599
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp -3599
transform -1 0 8464 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp -3599
transform -1 0 6808 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp -3599
transform -1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp -3599
transform 1 0 7636 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp -3599
transform 1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp -3599
transform 1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1011_
timestamp -3599
transform 1 0 13064 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1012_
timestamp -3599
transform 1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp -3599
transform -1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp -3599
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp -3599
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp -3599
transform 1 0 14996 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp -3599
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp -3599
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp -3599
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp -3599
transform -1 0 21804 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp -3599
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp -3599
transform -1 0 24104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp -3599
transform -1 0 24104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp -3599
transform 1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp -3599
transform 1 0 14720 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp -3599
transform 1 0 14168 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp -3599
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp -3599
transform 1 0 12788 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp -3599
transform -1 0 10028 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp -3599
transform -1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp -3599
transform -1 0 8924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp -3599
transform -1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp -3599
transform -1 0 9200 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp -3599
transform -1 0 10672 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp -3599
transform -1 0 10212 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp -3599
transform -1 0 11040 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp -3599
transform -1 0 11316 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp -3599
transform -1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp -3599
transform -1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp -3599
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp -3599
transform -1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp -3599
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp -3599
transform -1 0 21528 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp -3599
transform -1 0 21344 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp -3599
transform 1 0 19412 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1046_
timestamp -3599
transform 1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1047_
timestamp -3599
transform -1 0 14720 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1048_
timestamp -3599
transform -1 0 8556 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp -3599
transform 1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp -3599
transform -1 0 6532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp -3599
transform 1 0 5888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp -3599
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp -3599
transform -1 0 6256 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp -3599
transform -1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp -3599
transform 1 0 8188 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp -3599
transform -1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp -3599
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp -3599
transform -1 0 8188 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp -3599
transform 1 0 23368 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1060_
timestamp -3599
transform -1 0 9568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1061_
timestamp -3599
transform -1 0 13432 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1062_
timestamp -3599
transform 1 0 12880 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1063_
timestamp -3599
transform -1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1064_
timestamp -3599
transform -1 0 9936 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1065_
timestamp -3599
transform 1 0 11408 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1066_
timestamp -3599
transform 1 0 10120 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1067_
timestamp -3599
transform -1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1068_
timestamp -3599
transform 1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp -3599
transform -1 0 11040 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1070_
timestamp -3599
transform -1 0 10120 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1071_
timestamp -3599
transform -1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1072_
timestamp -3599
transform -1 0 11408 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1073_
timestamp -3599
transform -1 0 13248 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1074_
timestamp -3599
transform -1 0 13616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1075_
timestamp -3599
transform 1 0 9108 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp -3599
transform 1 0 10764 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1077_
timestamp -3599
transform 1 0 21988 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1078_
timestamp -3599
transform -1 0 22908 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1079_
timestamp -3599
transform 1 0 21528 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1080_
timestamp -3599
transform -1 0 22816 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp -3599
transform -1 0 19044 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1082_
timestamp -3599
transform -1 0 21528 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1083_
timestamp -3599
transform -1 0 21528 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1084_
timestamp -3599
transform 1 0 19136 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1085_
timestamp -3599
transform -1 0 19136 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1086_
timestamp -3599
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1087_
timestamp -3599
transform 1 0 15272 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp -3599
transform 1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1089_
timestamp -3599
transform 1 0 10120 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _1090_
timestamp -3599
transform 1 0 10120 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1091_
timestamp -3599
transform -1 0 10948 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp -3599
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1093_
timestamp -3599
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1094_
timestamp -3599
transform 1 0 11776 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp -3599
transform -1 0 13340 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1096_
timestamp -3599
transform 1 0 9844 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1097_
timestamp -3599
transform 1 0 11040 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1098_
timestamp -3599
transform 1 0 12144 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1099_
timestamp -3599
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1100_
timestamp -3599
transform 1 0 13340 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1101_
timestamp -3599
transform 1 0 12696 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1102_
timestamp -3599
transform 1 0 12604 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _1103_
timestamp -3599
transform 1 0 13432 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1104_
timestamp -3599
transform -1 0 12328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1105_
timestamp -3599
transform -1 0 13432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1106_
timestamp -3599
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1107_
timestamp -3599
transform 1 0 12420 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1108_
timestamp -3599
transform -1 0 18308 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1109_
timestamp -3599
transform -1 0 14628 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1110_
timestamp -3599
transform -1 0 14996 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1111_
timestamp -3599
transform -1 0 18768 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1112_
timestamp -3599
transform 1 0 16652 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1113_
timestamp -3599
transform -1 0 16376 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1114_
timestamp -3599
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1115_
timestamp -3599
transform 1 0 14260 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1116_
timestamp -3599
transform 1 0 17480 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1117_
timestamp -3599
transform -1 0 17664 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1118_
timestamp -3599
transform -1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1119_
timestamp -3599
transform -1 0 15364 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp -3599
transform 1 0 15640 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1121_
timestamp -3599
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1122_
timestamp -3599
transform -1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1123_
timestamp -3599
transform -1 0 15916 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1124_
timestamp -3599
transform -1 0 23368 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp -3599
transform -1 0 21712 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1126_
timestamp -3599
transform -1 0 21712 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1127_
timestamp -3599
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1128_
timestamp -3599
transform 1 0 19688 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1129_
timestamp -3599
transform 1 0 20700 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1130_
timestamp -3599
transform 1 0 8096 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp -3599
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1132_
timestamp -3599
transform 1 0 10488 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1133_
timestamp -3599
transform 1 0 11040 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1134_
timestamp -3599
transform -1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1135_
timestamp -3599
transform -1 0 6808 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1136_
timestamp -3599
transform 1 0 6164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp -3599
transform 1 0 6716 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1138_
timestamp -3599
transform -1 0 13984 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_4  _1139_
timestamp -3599
transform 1 0 14168 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1140_
timestamp -3599
transform -1 0 19044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp -3599
transform 1 0 19044 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1142_
timestamp -3599
transform -1 0 19320 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp -3599
transform -1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp -3599
transform -1 0 20516 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1145_
timestamp -3599
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1146_
timestamp -3599
transform -1 0 21528 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1147_
timestamp -3599
transform 1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp -3599
transform 1 0 21620 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1149_
timestamp -3599
transform 1 0 22264 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1150_
timestamp -3599
transform -1 0 22816 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1151_
timestamp -3599
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1152_
timestamp -3599
transform -1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1153_
timestamp -3599
transform -1 0 21344 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1154_
timestamp -3599
transform 1 0 20332 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1155_
timestamp -3599
transform -1 0 19964 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1156_
timestamp -3599
transform 1 0 16744 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1157_
timestamp -3599
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1158_
timestamp -3599
transform -1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1159_
timestamp -3599
transform 1 0 16008 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1160_
timestamp -3599
transform -1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1161_
timestamp -3599
transform -1 0 17572 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1162_
timestamp -3599
transform -1 0 17572 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1163_
timestamp -3599
transform 1 0 17296 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1164_
timestamp -3599
transform -1 0 18768 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1165_
timestamp -3599
transform 1 0 6072 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1166_
timestamp -3599
transform -1 0 7636 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1167_
timestamp -3599
transform 1 0 2760 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1168_
timestamp -3599
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp -3599
transform -1 0 7636 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1170_
timestamp -3599
transform 1 0 5796 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1171_
timestamp -3599
transform -1 0 5336 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1172_
timestamp -3599
transform 1 0 5612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1173_
timestamp -3599
transform -1 0 7268 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp -3599
transform 1 0 2576 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp -3599
transform -1 0 3680 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp -3599
transform 1 0 3036 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1177_
timestamp -3599
transform -1 0 4416 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1178_
timestamp -3599
transform -1 0 5152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp -3599
transform -1 0 4140 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1180_
timestamp -3599
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1181_
timestamp -3599
transform 1 0 4968 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1182_
timestamp -3599
transform -1 0 4876 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1183_
timestamp -3599
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1184_
timestamp -3599
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1185_
timestamp -3599
transform 1 0 5244 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1186_
timestamp -3599
transform -1 0 2760 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1187_
timestamp -3599
transform 1 0 4416 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp -3599
transform -1 0 3220 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1189_
timestamp -3599
transform -1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1190_
timestamp -3599
transform -1 0 5796 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1191_
timestamp -3599
transform -1 0 5888 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1192_
timestamp -3599
transform 1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1193_
timestamp -3599
transform 1 0 5060 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1194_
timestamp -3599
transform 1 0 7268 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1195_
timestamp -3599
transform 1 0 8096 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1196_
timestamp -3599
transform 1 0 9660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp -3599
transform -1 0 10488 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp -3599
transform -1 0 11040 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1199_
timestamp -3599
transform 1 0 10580 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1200_
timestamp -3599
transform -1 0 14628 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp -3599
transform -1 0 11408 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1202_
timestamp -3599
transform 1 0 11408 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1203_
timestamp -3599
transform -1 0 12420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1204_
timestamp -3599
transform 1 0 18492 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1205_
timestamp -3599
transform -1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp -3599
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1207_
timestamp -3599
transform -1 0 19412 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1208_
timestamp -3599
transform 1 0 16744 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp -3599
transform 1 0 18032 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1210_
timestamp -3599
transform -1 0 17296 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1211_
timestamp -3599
transform -1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1212_
timestamp -3599
transform 1 0 18216 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1213_
timestamp -3599
transform 1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1214_
timestamp -3599
transform -1 0 18124 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _1215_
timestamp -3599
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1216_
timestamp -3599
transform -1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1217_
timestamp -3599
transform 1 0 21804 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1218_
timestamp -3599
transform -1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp -3599
transform 1 0 20700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1220_
timestamp -3599
transform 1 0 21712 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1221_
timestamp -3599
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1222_
timestamp -3599
transform 1 0 22264 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1223_
timestamp -3599
transform 1 0 21712 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1224_
timestamp -3599
transform -1 0 22448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1225_
timestamp -3599
transform 1 0 22632 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1226_
timestamp -3599
transform -1 0 21712 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1227_
timestamp -3599
transform 1 0 21988 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1228_
timestamp -3599
transform 1 0 21988 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1229_
timestamp -3599
transform 1 0 23184 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1230_
timestamp -3599
transform -1 0 18216 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1231_
timestamp -3599
transform -1 0 18032 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp -3599
transform 1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1233_
timestamp -3599
transform -1 0 18400 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1234_
timestamp -3599
transform 1 0 18492 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1235_
timestamp -3599
transform 1 0 19780 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1236_
timestamp -3599
transform -1 0 17572 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1237_
timestamp -3599
transform 1 0 15640 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp -3599
transform 1 0 18032 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1239_
timestamp -3599
transform -1 0 19780 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp -3599
transform 1 0 15456 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1241_
timestamp -3599
transform 1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1242_
timestamp -3599
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1243_
timestamp -3599
transform -1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1244_
timestamp -3599
transform -1 0 10580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1245_
timestamp -3599
transform -1 0 10580 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1246_
timestamp -3599
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1247_
timestamp -3599
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1248_
timestamp -3599
transform -1 0 9384 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1249_
timestamp -3599
transform 1 0 7084 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1250_
timestamp -3599
transform 1 0 13064 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1251_
timestamp -3599
transform -1 0 13064 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1252_
timestamp -3599
transform 1 0 12696 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1253_
timestamp -3599
transform 1 0 10764 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1254_
timestamp -3599
transform 1 0 11776 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1255_
timestamp -3599
transform -1 0 9108 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1256_
timestamp -3599
transform 1 0 6532 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp -3599
transform -1 0 3680 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp -3599
transform 1 0 3312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_1  _1259_
timestamp -3599
transform 1 0 3772 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1260_
timestamp -3599
transform -1 0 4324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1261_
timestamp -3599
transform 1 0 4508 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1262_
timestamp -3599
transform 1 0 4692 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1263_
timestamp -3599
transform 1 0 3772 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1264_
timestamp -3599
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1265_
timestamp -3599
transform 1 0 1932 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1266_
timestamp -3599
transform 1 0 2208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1267_
timestamp -3599
transform -1 0 5244 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp -3599
transform -1 0 3680 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1269_
timestamp -3599
transform -1 0 4416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1270_
timestamp -3599
transform 1 0 4876 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1271_
timestamp -3599
transform 1 0 4140 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1272_
timestamp -3599
transform -1 0 4048 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1273_
timestamp -3599
transform -1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1274_
timestamp -3599
transform 1 0 2484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1275_
timestamp -3599
transform 1 0 2484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp -3599
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1277_
timestamp -3599
transform 1 0 1380 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1278_
timestamp -3599
transform 1 0 1840 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1279_
timestamp -3599
transform -1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1280_
timestamp -3599
transform 1 0 2300 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _1281_
timestamp -3599
transform 1 0 5428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp -3599
transform -1 0 5152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp -3599
transform 1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1284_
timestamp -3599
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1285_
timestamp -3599
transform -1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1286_
timestamp -3599
transform 1 0 4048 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1287_
timestamp -3599
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1288_
timestamp -3599
transform 1 0 4232 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1289_
timestamp -3599
transform 1 0 4692 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1290_
timestamp -3599
transform -1 0 3956 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1291_
timestamp -3599
transform 1 0 2484 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1292_
timestamp -3599
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1293_
timestamp -3599
transform 1 0 6624 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21bai_1  _1294_
timestamp -3599
transform 1 0 6624 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1295_
timestamp -3599
transform 1 0 6900 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1296_
timestamp -3599
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp -3599
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1298_
timestamp -3599
transform -1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1299_
timestamp -3599
transform 1 0 16928 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1300_
timestamp -3599
transform -1 0 17296 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1301_
timestamp -3599
transform 1 0 15180 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1302_
timestamp -3599
transform 1 0 17664 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1303_
timestamp -3599
transform -1 0 19688 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1304_
timestamp -3599
transform 1 0 16928 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1305_
timestamp -3599
transform 1 0 17204 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1306_
timestamp -3599
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1307_
timestamp -3599
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1308_
timestamp -3599
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1309_
timestamp -3599
transform -1 0 21528 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1310_
timestamp -3599
transform 1 0 21528 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1311_
timestamp -3599
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1312_
timestamp -3599
transform 1 0 20240 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1313_
timestamp -3599
transform 1 0 20884 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1314_
timestamp -3599
transform 1 0 23000 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp -3599
transform 1 0 24380 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1316_
timestamp -3599
transform 1 0 21896 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1317_
timestamp -3599
transform 1 0 27508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1318_
timestamp -3599
transform 1 0 27416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1319_
timestamp -3599
transform -1 0 26864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1320_
timestamp -3599
transform 1 0 26956 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp -3599
transform -1 0 27600 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1322_
timestamp -3599
transform -1 0 28244 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp -3599
transform 1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1324_
timestamp -3599
transform 1 0 26220 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1325_
timestamp -3599
transform 1 0 27600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1326_
timestamp -3599
transform -1 0 27600 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp -3599
transform -1 0 26680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1328_
timestamp -3599
transform 1 0 26864 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1329_
timestamp -3599
transform 1 0 27140 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1330_
timestamp -3599
transform -1 0 27692 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1331_
timestamp -3599
transform 1 0 27232 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1332_
timestamp -3599
transform -1 0 28060 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1333_
timestamp -3599
transform -1 0 26036 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1334_
timestamp -3599
transform -1 0 24380 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1335_
timestamp -3599
transform 1 0 23552 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1336_
timestamp -3599
transform -1 0 24104 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1337_
timestamp -3599
transform 1 0 17848 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1338_
timestamp -3599
transform 1 0 16652 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1339_
timestamp -3599
transform 1 0 15180 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_1  _1340_
timestamp -3599
transform 1 0 14168 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1341_
timestamp -3599
transform -1 0 16376 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1342_
timestamp -3599
transform 1 0 17296 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1343_
timestamp -3599
transform 1 0 16744 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1344_
timestamp -3599
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1345_
timestamp -3599
transform -1 0 19044 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1346_
timestamp -3599
transform 1 0 16008 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1347_
timestamp -3599
transform 1 0 18492 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1348_
timestamp -3599
transform 1 0 13524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1349_
timestamp -3599
transform -1 0 13524 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1350_
timestamp -3599
transform -1 0 13708 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1351_
timestamp -3599
transform 1 0 10120 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1352_
timestamp -3599
transform -1 0 11408 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1353_
timestamp -3599
transform -1 0 9568 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1354_
timestamp -3599
transform 1 0 9292 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1355_
timestamp -3599
transform 1 0 9384 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1356_
timestamp -3599
transform 1 0 9568 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp -3599
transform 1 0 10580 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1358_
timestamp -3599
transform -1 0 11040 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1359_
timestamp -3599
transform 1 0 11132 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1360_
timestamp -3599
transform 1 0 13340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1361_
timestamp -3599
transform -1 0 19688 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1362_
timestamp -3599
transform -1 0 22908 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1363_
timestamp -3599
transform -1 0 23368 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1364_
timestamp -3599
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1365_
timestamp -3599
transform -1 0 22816 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1366_
timestamp -3599
transform 1 0 20884 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1367_
timestamp -3599
transform -1 0 20332 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1368_
timestamp -3599
transform 1 0 20056 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1369_
timestamp -3599
transform 1 0 18584 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1370_
timestamp -3599
transform 1 0 15916 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp -3599
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1372_
timestamp -3599
transform -1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp -3599
transform 1 0 12236 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1374_
timestamp -3599
transform 1 0 12880 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1375_
timestamp -3599
transform -1 0 13892 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1376_
timestamp -3599
transform -1 0 14168 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1377_
timestamp -3599
transform 1 0 12052 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1378_
timestamp -3599
transform 1 0 12696 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1379_
timestamp -3599
transform 1 0 11868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1380_
timestamp -3599
transform -1 0 13156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1381_
timestamp -3599
transform -1 0 14720 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1382_
timestamp -3599
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp -3599
transform 1 0 13616 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp -3599
transform -1 0 13524 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1385_
timestamp -3599
transform 1 0 13248 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1386_
timestamp -3599
transform -1 0 12880 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1387_
timestamp -3599
transform 1 0 13156 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1388_
timestamp -3599
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1389_
timestamp -3599
transform 1 0 12420 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1390_
timestamp -3599
transform 1 0 13524 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp -3599
transform 1 0 12604 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1392_
timestamp -3599
transform -1 0 11960 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp -3599
transform 1 0 12236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1394_
timestamp -3599
transform 1 0 12420 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1395_
timestamp -3599
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1396_
timestamp -3599
transform 1 0 12604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1397_
timestamp -3599
transform 1 0 16836 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1398_
timestamp -3599
transform -1 0 16560 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1399_
timestamp -3599
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp -3599
transform 1 0 15180 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1401_
timestamp -3599
transform -1 0 15180 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1402_
timestamp -3599
transform 1 0 14812 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1403_
timestamp -3599
transform 1 0 14628 0 1 26112
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _1404_
timestamp -3599
transform 1 0 23368 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1405_
timestamp -3599
transform -1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1406_
timestamp -3599
transform 1 0 22816 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1407_
timestamp -3599
transform 1 0 23184 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1408_
timestamp -3599
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1409_
timestamp -3599
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1410_
timestamp -3599
transform 1 0 20700 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1411_
timestamp -3599
transform 1 0 22540 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp -3599
transform -1 0 20700 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1413_
timestamp -3599
transform 1 0 19412 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1414_
timestamp -3599
transform -1 0 18216 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1415_
timestamp -3599
transform 1 0 18032 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1416_
timestamp -3599
transform 1 0 18492 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1417_
timestamp -3599
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp -3599
transform -1 0 16560 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1419_
timestamp -3599
transform 1 0 16192 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1420_
timestamp -3599
transform 1 0 17388 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1421_
timestamp -3599
transform -1 0 16376 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1422_
timestamp -3599
transform 1 0 14352 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1423_
timestamp -3599
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1424_
timestamp -3599
transform 1 0 12972 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1425_
timestamp -3599
transform -1 0 13892 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp -3599
transform 1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1427_
timestamp -3599
transform -1 0 11776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1428_
timestamp -3599
transform 1 0 10304 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1429_
timestamp -3599
transform 1 0 12512 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp -3599
transform 1 0 10948 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1431_
timestamp -3599
transform -1 0 12144 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1432_
timestamp -3599
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1433_
timestamp -3599
transform 1 0 13064 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1434_
timestamp -3599
transform 1 0 13524 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1435_
timestamp -3599
transform -1 0 14168 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1436_
timestamp -3599
transform -1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1437_
timestamp -3599
transform 1 0 14168 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1438_
timestamp -3599
transform -1 0 13984 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp -3599
transform 1 0 14720 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1440_
timestamp -3599
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1441_
timestamp -3599
transform -1 0 6716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1442_
timestamp -3599
transform -1 0 6532 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1443_
timestamp -3599
transform -1 0 6440 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1444_
timestamp -3599
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1445_
timestamp -3599
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1446_
timestamp -3599
transform 1 0 6348 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1447_
timestamp -3599
transform -1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1448_
timestamp -3599
transform -1 0 6808 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1449_
timestamp -3599
transform -1 0 5152 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1450_
timestamp -3599
transform -1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1451_
timestamp -3599
transform -1 0 5152 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1452_
timestamp -3599
transform -1 0 4692 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1453_
timestamp -3599
transform 1 0 4140 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp -3599
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1455_
timestamp -3599
transform -1 0 4600 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1456_
timestamp -3599
transform -1 0 5060 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1457_
timestamp -3599
transform 1 0 4232 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1458_
timestamp -3599
transform -1 0 4784 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1459_
timestamp -3599
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp -3599
transform -1 0 7176 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1461_
timestamp -3599
transform -1 0 6808 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1462_
timestamp -3599
transform -1 0 7176 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1463_
timestamp -3599
transform 1 0 7176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1464_
timestamp -3599
transform -1 0 8740 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp -3599
transform 1 0 7452 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1466_
timestamp -3599
transform -1 0 8280 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1467_
timestamp -3599
transform -1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp -3599
transform 1 0 9844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1469_
timestamp -3599
transform -1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1470_
timestamp -3599
transform 1 0 10948 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1471_
timestamp -3599
transform 1 0 10672 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1472_
timestamp -3599
transform 1 0 10672 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1473_
timestamp -3599
transform 1 0 13156 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1474_
timestamp -3599
transform -1 0 14168 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1475_
timestamp -3599
transform -1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1476_
timestamp -3599
transform 1 0 14444 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1477_
timestamp -3599
transform 1 0 14168 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1478_
timestamp -3599
transform -1 0 15180 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1479_
timestamp -3599
transform 1 0 15456 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1480_
timestamp -3599
transform 1 0 15272 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1481_
timestamp -3599
transform 1 0 15732 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp -3599
transform 1 0 17664 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1483_
timestamp -3599
transform 1 0 17204 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1484_
timestamp -3599
transform 1 0 17480 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1485_
timestamp -3599
transform 1 0 19136 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp -3599
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1487_
timestamp -3599
transform 1 0 19596 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1488_
timestamp -3599
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1489_
timestamp -3599
transform 1 0 18676 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1490_
timestamp -3599
transform 1 0 19504 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1491_
timestamp -3599
transform 1 0 19872 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1492_
timestamp -3599
transform 1 0 19596 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1493_
timestamp -3599
transform 1 0 20332 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1494_
timestamp -3599
transform 1 0 19320 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1495_
timestamp -3599
transform 1 0 14260 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1496_
timestamp -3599
transform -1 0 24012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1497_
timestamp -3599
transform -1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1498_
timestamp -3599
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _1499_
timestamp -3599
transform 1 0 22908 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1500_
timestamp -3599
transform -1 0 13248 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1501_
timestamp -3599
transform 1 0 9660 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1502_
timestamp -3599
transform 1 0 6992 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1503_
timestamp -3599
transform 1 0 7360 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1504_
timestamp -3599
transform -1 0 8924 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp -3599
transform 1 0 10304 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1506_
timestamp -3599
transform 1 0 10764 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1507_
timestamp -3599
transform 1 0 9292 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1508_
timestamp -3599
transform -1 0 10488 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1509_
timestamp -3599
transform -1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1510_
timestamp -3599
transform -1 0 13340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1511_
timestamp -3599
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1512_
timestamp -3599
transform 1 0 24104 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1513_
timestamp -3599
transform -1 0 25392 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1514_
timestamp -3599
transform -1 0 25024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1515_
timestamp -3599
transform -1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1516_
timestamp -3599
transform -1 0 21620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1517_
timestamp -3599
transform 1 0 18492 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp -3599
transform 1 0 17112 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1519_
timestamp -3599
transform 1 0 17756 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1520_
timestamp -3599
transform 1 0 14812 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1521_
timestamp -3599
transform 1 0 13248 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1522_
timestamp -3599
transform 1 0 14168 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1523_
timestamp -3599
transform 1 0 13340 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp -3599
transform -1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1525_
timestamp -3599
transform 1 0 13800 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp -3599
transform 1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1527_
timestamp -3599
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1528_
timestamp -3599
transform 1 0 9936 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp -3599
transform 1 0 10396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1530_
timestamp -3599
transform 1 0 10764 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1531_
timestamp -3599
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1532_
timestamp -3599
transform -1 0 11132 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o32ai_1  _1533_
timestamp -3599
transform 1 0 11500 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1534_
timestamp -3599
transform 1 0 11592 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1535_
timestamp -3599
transform 1 0 12144 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1536_
timestamp -3599
transform -1 0 12696 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1537_
timestamp -3599
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1538_
timestamp -3599
transform 1 0 11868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1539_
timestamp -3599
transform 1 0 10488 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1540_
timestamp -3599
transform 1 0 10856 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1541_
timestamp -3599
transform 1 0 12236 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1542_
timestamp -3599
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp -3599
transform -1 0 17296 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1544_
timestamp -3599
transform 1 0 18308 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp -3599
transform 1 0 14444 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1546_
timestamp -3599
transform -1 0 16744 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp -3599
transform -1 0 19596 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp -3599
transform 1 0 17572 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1549_
timestamp -3599
transform -1 0 17112 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1550_
timestamp -3599
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1551_
timestamp -3599
transform -1 0 15640 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1552_
timestamp -3599
transform 1 0 13800 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1553_
timestamp -3599
transform -1 0 16008 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1554_
timestamp -3599
transform -1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1555_
timestamp -3599
transform -1 0 17388 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1556_
timestamp -3599
transform 1 0 18492 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1557_
timestamp -3599
transform -1 0 18492 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1558_
timestamp -3599
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1559_
timestamp -3599
transform 1 0 9108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1560_
timestamp -3599
transform -1 0 9108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1561_
timestamp -3599
transform 1 0 9200 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp -3599
transform 1 0 9016 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1563_
timestamp -3599
transform -1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1564_
timestamp -3599
transform -1 0 23000 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1565_
timestamp -3599
transform 1 0 22632 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1566_
timestamp -3599
transform 1 0 23276 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1567_
timestamp -3599
transform -1 0 22448 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1568_
timestamp -3599
transform -1 0 20700 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1569_
timestamp -3599
transform 1 0 17204 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1570_
timestamp -3599
transform 1 0 18400 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1571_
timestamp -3599
transform 1 0 17848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1572_
timestamp -3599
transform 1 0 14904 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1573_
timestamp -3599
transform -1 0 13340 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1574_
timestamp -3599
transform 1 0 14168 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1575_
timestamp -3599
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1576_
timestamp -3599
transform -1 0 12144 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1577_
timestamp -3599
transform 1 0 11500 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1578_
timestamp -3599
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1579_
timestamp -3599
transform -1 0 12236 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1580_
timestamp -3599
transform -1 0 10764 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1581_
timestamp -3599
transform 1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp -3599
transform -1 0 8188 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1583_
timestamp -3599
transform 1 0 5612 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1584_
timestamp -3599
transform 1 0 6992 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1585_
timestamp -3599
transform 1 0 5244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1586_
timestamp -3599
transform 1 0 5336 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1587_
timestamp -3599
transform 1 0 7544 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1588_
timestamp -3599
transform 1 0 6164 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1589_
timestamp -3599
transform -1 0 7176 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1590_
timestamp -3599
transform 1 0 5888 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1591_
timestamp -3599
transform 1 0 8188 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1592_
timestamp -3599
transform 1 0 5428 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1593_
timestamp -3599
transform 1 0 5796 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1594_
timestamp -3599
transform 1 0 6440 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1595_
timestamp -3599
transform 1 0 7360 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1596_
timestamp -3599
transform 1 0 7728 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1597_
timestamp -3599
transform -1 0 9660 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1598_
timestamp -3599
transform 1 0 19688 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp -3599
transform 1 0 20976 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1600_
timestamp -3599
transform -1 0 21252 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1601_
timestamp -3599
transform 1 0 14996 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1602_
timestamp -3599
transform -1 0 20700 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1603_
timestamp -3599
transform 1 0 21620 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp -3599
transform -1 0 20240 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1605_
timestamp -3599
transform -1 0 14812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1606_
timestamp -3599
transform 1 0 15640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _1607_
timestamp -3599
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1608_
timestamp -3599
transform 1 0 18400 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp -3599
transform 1 0 18676 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1610_
timestamp -3599
transform -1 0 20976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1611_
timestamp -3599
transform -1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1612_
timestamp -3599
transform 1 0 19780 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1613_
timestamp -3599
transform 1 0 10396 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1614_
timestamp -3599
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1615_
timestamp -3599
transform 1 0 16744 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1616_
timestamp -3599
transform -1 0 25024 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1617_
timestamp -3599
transform -1 0 24656 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1618_
timestamp -3599
transform 1 0 23092 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1619_
timestamp -3599
transform 1 0 23736 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1620_
timestamp -3599
transform 1 0 20056 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1621_
timestamp -3599
transform -1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp -3599
transform 1 0 19320 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp -3599
transform -1 0 17480 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1624_
timestamp -3599
transform 1 0 14444 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp -3599
transform 1 0 10028 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1626_
timestamp -3599
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1627_
timestamp -3599
transform 1 0 10672 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1628_
timestamp -3599
transform 1 0 9936 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1629_
timestamp -3599
transform 1 0 10028 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1630_
timestamp -3599
transform 1 0 10948 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1631_
timestamp -3599
transform 1 0 10304 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1632_
timestamp -3599
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1633_
timestamp -3599
transform 1 0 9660 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp -3599
transform 1 0 10488 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_2  _1635_
timestamp -3599
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp -3599
transform -1 0 10396 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp -3599
transform 1 0 8740 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1638_
timestamp -3599
transform 1 0 9292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1639_
timestamp -3599
transform 1 0 13524 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp -3599
transform -1 0 11224 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp -3599
transform 1 0 7452 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1642_
timestamp -3599
transform -1 0 8004 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1643_
timestamp -3599
transform -1 0 13248 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1644_
timestamp -3599
transform -1 0 12328 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1645_
timestamp -3599
transform 1 0 8188 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1646_
timestamp -3599
transform -1 0 11132 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _1647_
timestamp -3599
transform -1 0 12788 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1648_
timestamp -3599
transform 1 0 7360 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1649_
timestamp -3599
transform 1 0 8188 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1650_
timestamp -3599
transform 1 0 8924 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1651_
timestamp -3599
transform -1 0 9660 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1652_
timestamp -3599
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1653_
timestamp -3599
transform -1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp -3599
transform 1 0 17664 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1655_
timestamp -3599
transform 1 0 14628 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1656_
timestamp -3599
transform -1 0 19044 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _1657_
timestamp -3599
transform 1 0 18308 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1658_
timestamp -3599
transform -1 0 18308 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1659_
timestamp -3599
transform 1 0 16652 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1660_
timestamp -3599
transform 1 0 17296 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1661_
timestamp -3599
transform -1 0 16560 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1662_
timestamp -3599
transform -1 0 17112 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1663_
timestamp -3599
transform 1 0 14168 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1664_
timestamp -3599
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1665_
timestamp -3599
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1666_
timestamp -3599
transform 1 0 15272 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1667_
timestamp -3599
transform 1 0 16376 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1668_
timestamp -3599
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _1669_
timestamp -3599
transform -1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1670_
timestamp -3599
transform 1 0 17848 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1671_
timestamp -3599
transform 1 0 19228 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1672_
timestamp -3599
transform 1 0 20884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1673_
timestamp -3599
transform 1 0 21620 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp -3599
transform 1 0 20884 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp -3599
transform 1 0 18768 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1676_
timestamp -3599
transform 1 0 15180 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1677_
timestamp -3599
transform 1 0 19044 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1678_
timestamp -3599
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1679_
timestamp -3599
transform 1 0 20976 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1680_
timestamp -3599
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1681_
timestamp -3599
transform 1 0 8096 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1682_
timestamp -3599
transform 1 0 8740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1683_
timestamp -3599
transform -1 0 8648 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1684_
timestamp -3599
transform 1 0 5336 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1685_
timestamp -3599
transform -1 0 6992 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1686_
timestamp -3599
transform -1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1687_
timestamp -3599
transform -1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1688_
timestamp -3599
transform -1 0 6624 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1689_
timestamp -3599
transform 1 0 5612 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1690_
timestamp -3599
transform 1 0 6348 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1691_
timestamp -3599
transform 1 0 7820 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp -3599
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1693_
timestamp -3599
transform 1 0 6716 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1694_
timestamp -3599
transform 1 0 20240 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1695_
timestamp -3599
transform -1 0 23920 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1696_
timestamp -3599
transform 1 0 23368 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1697_
timestamp -3599
transform 1 0 22080 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1698_
timestamp -3599
transform -1 0 23736 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp -3599
transform -1 0 20792 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1700_
timestamp -3599
transform 1 0 18032 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1701_
timestamp -3599
transform -1 0 18032 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1702_
timestamp -3599
transform 1 0 17296 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1703_
timestamp -3599
transform -1 0 15916 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1704_
timestamp -3599
transform -1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1705_
timestamp -3599
transform 1 0 8740 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1706_
timestamp -3599
transform 1 0 8280 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1707_
timestamp -3599
transform -1 0 8740 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp -3599
transform -1 0 9476 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1709_
timestamp -3599
transform 1 0 7728 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1710_
timestamp -3599
transform -1 0 9384 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1711_
timestamp -3599
transform 1 0 8372 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1712_
timestamp -3599
transform 1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1713_
timestamp -3599
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1714_
timestamp -3599
transform 1 0 7452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1715_
timestamp -3599
transform -1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1716_
timestamp -3599
transform -1 0 8096 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1717_
timestamp -3599
transform -1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1718_
timestamp -3599
transform 1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1719_
timestamp -3599
transform 1 0 8740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1720_
timestamp -3599
transform -1 0 8096 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1721_
timestamp -3599
transform -1 0 8740 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1722_
timestamp -3599
transform 1 0 7544 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1723_
timestamp -3599
transform 1 0 7360 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1724_
timestamp -3599
transform 1 0 6532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1725_
timestamp -3599
transform 1 0 6440 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1726_
timestamp -3599
transform 1 0 7728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1727_
timestamp -3599
transform -1 0 8004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1728_
timestamp -3599
transform 1 0 14628 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1729_
timestamp -3599
transform -1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1730_
timestamp -3599
transform 1 0 19964 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1731_
timestamp -3599
transform 1 0 19688 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1732_
timestamp -3599
transform 1 0 19412 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1733_
timestamp -3599
transform -1 0 20700 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1734_
timestamp -3599
transform 1 0 25760 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1735_
timestamp -3599
transform -1 0 27600 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1736_
timestamp -3599
transform 1 0 27968 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1737_
timestamp -3599
transform 1 0 28060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1738_
timestamp -3599
transform -1 0 27600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1739_
timestamp -3599
transform -1 0 28060 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1740_
timestamp -3599
transform -1 0 26128 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1741_
timestamp -3599
transform -1 0 25668 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1742_
timestamp -3599
transform -1 0 27600 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1743_
timestamp -3599
transform 1 0 27140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1744_
timestamp -3599
transform 1 0 27140 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1745_
timestamp -3599
transform -1 0 28704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1746_
timestamp -3599
transform 1 0 26956 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1747_
timestamp -3599
transform 1 0 26956 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1748_
timestamp -3599
transform -1 0 25944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1749_
timestamp -3599
transform -1 0 25852 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1750_
timestamp -3599
transform 1 0 25208 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1751_
timestamp -3599
transform 1 0 25116 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1752_
timestamp -3599
transform -1 0 27600 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1753_
timestamp -3599
transform 1 0 27048 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp -3599
transform 1 0 27324 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1755_
timestamp -3599
transform 1 0 27784 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1756_
timestamp -3599
transform 1 0 27324 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1757_
timestamp -3599
transform 1 0 26772 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1758_
timestamp -3599
transform -1 0 25668 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1759_
timestamp -3599
transform 1 0 25484 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1760_
timestamp -3599
transform -1 0 26404 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1761_
timestamp -3599
transform 1 0 24380 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1762_
timestamp -3599
transform -1 0 27508 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1763_
timestamp -3599
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1764_
timestamp -3599
transform 1 0 27416 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1765_
timestamp -3599
transform -1 0 28336 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1766_
timestamp -3599
transform 1 0 27600 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1767_
timestamp -3599
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1768_
timestamp -3599
transform -1 0 26864 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1769_
timestamp -3599
transform 1 0 27140 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1770_
timestamp -3599
transform 1 0 27600 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1771_
timestamp -3599
transform 1 0 27140 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1772_
timestamp -3599
transform 1 0 26772 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1773_
timestamp -3599
transform -1 0 26036 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1774_
timestamp -3599
transform 1 0 26956 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1775_
timestamp -3599
transform -1 0 25852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1776_
timestamp -3599
transform -1 0 25392 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1777_
timestamp -3599
transform -1 0 24656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1778_
timestamp -3599
transform -1 0 24288 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1779_
timestamp -3599
transform 1 0 23276 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1780_
timestamp -3599
transform -1 0 23552 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1781_
timestamp -3599
transform 1 0 24012 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1782_
timestamp -3599
transform 1 0 23644 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1783_
timestamp -3599
transform 1 0 23184 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1784_
timestamp -3599
transform -1 0 23460 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_1  _1785_
timestamp -3599
transform -1 0 24932 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1786_
timestamp -3599
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1787_
timestamp -3599
transform -1 0 22080 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1788_
timestamp -3599
transform -1 0 24288 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp -3599
transform -1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1790_
timestamp -3599
transform 1 0 17664 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1791_
timestamp -3599
transform -1 0 20240 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1792_
timestamp -3599
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp -3599
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1794_
timestamp -3599
transform -1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1795_
timestamp -3599
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp -3599
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1797_
timestamp -3599
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1798_
timestamp -3599
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1799_
timestamp -3599
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1800_
timestamp -3599
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1801_
timestamp -3599
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1802_
timestamp -3599
transform 1 0 2300 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1803_
timestamp -3599
transform -1 0 4232 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1804_
timestamp -3599
transform 1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1805_
timestamp -3599
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1806_
timestamp -3599
transform -1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1807_
timestamp -3599
transform 1 0 14260 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1808_
timestamp -3599
transform 1 0 6808 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1809_
timestamp -3599
transform 1 0 16192 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp -3599
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1811_
timestamp -3599
transform -1 0 16928 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp -3599
transform -1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1813_
timestamp -3599
transform -1 0 24656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1814_
timestamp -3599
transform -1 0 25024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1815_
timestamp -3599
transform -1 0 24656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1816_
timestamp -3599
transform -1 0 24288 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1817_
timestamp -3599
transform -1 0 25208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1818_
timestamp -3599
transform -1 0 26404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1819_
timestamp -3599
transform 1 0 27232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1820_
timestamp -3599
transform -1 0 29164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp -3599
transform -1 0 28980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1822_
timestamp -3599
transform -1 0 27508 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1823_
timestamp -3599
transform -1 0 26496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1824_
timestamp -3599
transform -1 0 28980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1825_
timestamp -3599
transform -1 0 29072 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1826_
timestamp -3599
transform -1 0 29072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1827_
timestamp -3599
transform -1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1828_
timestamp -3599
transform 1 0 26128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1829_
timestamp -3599
transform 1 0 26220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp -3599
transform -1 0 28796 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1831_
timestamp -3599
transform -1 0 28980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1832_
timestamp -3599
transform -1 0 29072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1833_
timestamp -3599
transform 1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1834_
timestamp -3599
transform 1 0 26036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1835_
timestamp -3599
transform -1 0 27232 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1836_
timestamp -3599
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp -3599
transform -1 0 29072 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1838_
timestamp -3599
transform -1 0 29072 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1839_
timestamp -3599
transform 1 0 26220 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1840_
timestamp -3599
transform -1 0 28980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1841_
timestamp -3599
transform -1 0 29072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1842_
timestamp -3599
transform -1 0 26312 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1843_
timestamp -3599
transform -1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp -3599
transform -1 0 26864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1845_
timestamp -3599
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1846_
timestamp -3599
transform 1 0 22540 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp -3599
transform -1 0 24932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1848_
timestamp -3599
transform -1 0 25392 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1849_
timestamp -3599
transform 1 0 22356 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1850_
timestamp -3599
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1851_
timestamp -3599
transform -1 0 23000 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1852_
timestamp -3599
transform 1 0 24472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1853_
timestamp -3599
transform -1 0 25392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1854_
timestamp -3599
transform -1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1855_
timestamp -3599
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1856_
timestamp -3599
transform -1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1857_
timestamp -3599
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1858_
timestamp -3599
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1859_
timestamp -3599
transform -1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1860_
timestamp -3599
transform 1 0 11960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1861_
timestamp -3599
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1862_
timestamp -3599
transform -1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1863_
timestamp -3599
transform -1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1864_
timestamp -3599
transform -1 0 15916 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1865_
timestamp -3599
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1866_
timestamp -3599
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1867_
timestamp -3599
transform 1 0 5336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1868_
timestamp -3599
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1869_
timestamp -3599
transform -1 0 3404 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1870_
timestamp -3599
transform 1 0 4692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1871_
timestamp -3599
transform 1 0 5796 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1872_
timestamp -3599
transform -1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1873_
timestamp -3599
transform -1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1874_
timestamp -3599
transform 1 0 11132 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1875_
timestamp -3599
transform 1 0 12328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1876_
timestamp -3599
transform 1 0 13616 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1877_
timestamp -3599
transform -1 0 15824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1878_
timestamp -3599
transform 1 0 16928 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1879_
timestamp -3599
transform 1 0 18768 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp -3599
transform -1 0 21344 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1881_
timestamp -3599
transform 1 0 21160 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1882_
timestamp -3599
transform 1 0 22172 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1883_
timestamp -3599
transform -1 0 21620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1884_
timestamp -3599
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1885_
timestamp -3599
transform 1 0 22448 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1886_
timestamp -3599
transform -1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _1887_
timestamp -3599
transform 1 0 22540 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1888_
timestamp -3599
transform 1 0 23644 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1889_
timestamp -3599
transform 1 0 20608 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1890_
timestamp -3599
transform 1 0 22816 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1891_
timestamp -3599
transform 1 0 18584 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1892_
timestamp -3599
transform 1 0 16652 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1893_
timestamp -3599
transform -1 0 21068 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1894_
timestamp -3599
transform 1 0 14444 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1895_
timestamp -3599
transform 1 0 6900 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1896_
timestamp -3599
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1897_
timestamp -3599
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1898_
timestamp -3599
transform 1 0 4140 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1899_
timestamp -3599
transform 1 0 3956 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1900_
timestamp -3599
transform 1 0 1380 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1901_
timestamp -3599
transform 1 0 1380 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1902_
timestamp -3599
transform 1 0 2392 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1903_
timestamp -3599
transform 1 0 1656 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1904_
timestamp -3599
transform 1 0 1380 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1905_
timestamp -3599
transform 1 0 2852 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1906_
timestamp -3599
transform 1 0 3496 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1907_
timestamp -3599
transform 1 0 6348 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1908_
timestamp -3599
transform 1 0 11776 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1909_
timestamp -3599
transform 1 0 13248 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1910_
timestamp -3599
transform 1 0 5980 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1911_
timestamp -3599
transform 1 0 15180 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1912_
timestamp -3599
transform -1 0 21344 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1913_
timestamp -3599
transform 1 0 14996 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1914_
timestamp -3599
transform 1 0 19688 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1915_
timestamp -3599
transform 1 0 23000 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1916_
timestamp -3599
transform 1 0 22908 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1917_
timestamp -3599
transform 1 0 23276 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1918_
timestamp -3599
transform -1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1919_
timestamp -3599
transform 1 0 23644 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1920_
timestamp -3599
transform 1 0 25024 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1921_
timestamp -3599
transform 1 0 26956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1922_
timestamp -3599
transform 1 0 27600 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1923_
timestamp -3599
transform 1 0 27600 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1924_
timestamp -3599
transform 1 0 25392 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1925_
timestamp -3599
transform 1 0 24656 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1926_
timestamp -3599
transform 1 0 27600 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1927_
timestamp -3599
transform 1 0 27600 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1928_
timestamp -3599
transform 1 0 27600 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1929_
timestamp -3599
transform 1 0 24840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1930_
timestamp -3599
transform 1 0 25116 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1931_
timestamp -3599
transform 1 0 25208 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1932_
timestamp -3599
transform 1 0 27416 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1933_
timestamp -3599
transform 1 0 27600 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1934_
timestamp -3599
transform 1 0 27600 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1935_
timestamp -3599
transform 1 0 24932 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1936_
timestamp -3599
transform 1 0 25024 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1937_
timestamp -3599
transform 1 0 25024 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1938_
timestamp -3599
transform 1 0 27508 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1939_
timestamp -3599
transform 1 0 27600 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1940_
timestamp -3599
transform 1 0 27600 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1941_
timestamp -3599
transform 1 0 25392 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1942_
timestamp -3599
transform 1 0 27600 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1943_
timestamp -3599
transform 1 0 27600 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1944_
timestamp -3599
transform 1 0 24932 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1945_
timestamp -3599
transform 1 0 27048 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1946_
timestamp -3599
transform 1 0 24748 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1947_
timestamp -3599
transform 1 0 22172 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1948_
timestamp -3599
transform -1 0 23920 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1949_
timestamp -3599
transform -1 0 25300 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1950_
timestamp -3599
transform -1 0 25944 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1951_
timestamp -3599
transform 1 0 21804 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1952_
timestamp -3599
transform 1 0 21804 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1953_
timestamp -3599
transform 1 0 20884 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1954_
timestamp -3599
transform 1 0 23460 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1955_
timestamp -3599
transform 1 0 23276 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1956_
timestamp -3599
transform 1 0 20700 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1957_
timestamp -3599
transform 1 0 19412 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1958_
timestamp -3599
transform -1 0 20332 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1959_
timestamp -3599
transform -1 0 18492 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1960_
timestamp -3599
transform 1 0 14352 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1961_
timestamp -3599
transform 1 0 12972 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1962_
timestamp -3599
transform 1 0 10948 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1963_
timestamp -3599
transform 1 0 8924 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1964_
timestamp -3599
transform -1 0 16008 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1965_
timestamp -3599
transform 1 0 14628 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1966_
timestamp -3599
transform 1 0 14536 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1967_
timestamp -3599
transform 1 0 4232 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1968_
timestamp -3599
transform 1 0 6992 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1969_
timestamp -3599
transform 1 0 4416 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1970_
timestamp -3599
transform 1 0 2760 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1971_
timestamp -3599
transform 1 0 1840 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1972_
timestamp -3599
transform 1 0 3680 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1973_
timestamp -3599
transform 1 0 4784 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1974_
timestamp -3599
transform 1 0 7820 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1975_
timestamp -3599
transform 1 0 7728 0 -1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1976_
timestamp -3599
transform 1 0 10120 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1977_
timestamp -3599
transform 1 0 11316 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1978_
timestamp -3599
transform 1 0 12604 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1979_
timestamp -3599
transform 1 0 14444 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1980_
timestamp -3599
transform -1 0 18584 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1981_
timestamp -3599
transform 1 0 17756 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1982_
timestamp -3599
transform 1 0 19964 0 1 28288
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1983_
timestamp -3599
transform 1 0 20148 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1984_
timestamp -3599
transform -1 0 23644 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1985_
timestamp -3599
transform 1 0 19872 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1986_
timestamp -3599
transform 1 0 22724 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1987_
timestamp -3599
transform 1 0 21436 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1988_
timestamp -3599
transform 1 0 14260 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp -3599
transform -1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3599
transform 1 0 15364 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp -3599
transform 1 0 6992 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp -3599
transform -1 0 13340 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp -3599
transform -1 0 8740 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp -3599
transform 1 0 10028 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp -3599
transform 1 0 21804 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp -3599
transform 1 0 24380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp -3599
transform -1 0 23276 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp -3599
transform 1 0 23644 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_8  clkload0
timestamp -3599
transform 1 0 7268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload1
timestamp -3599
transform 1 0 11316 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload2
timestamp -3599
transform 1 0 6900 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_12  clkload3
timestamp -3599
transform 1 0 10028 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload4
timestamp -3599
transform 1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload5
timestamp -3599
transform 1 0 23644 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp -3599
transform 1 0 20792 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20
timestamp -3599
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43
timestamp -3599
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp -3599
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp -3599
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp -3599
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp -3599
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp -3599
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp -3599
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp -3599
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp -3599
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp -3599
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_119
timestamp -3599
transform 1 0 12052 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp -3599
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp -3599
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp -3599
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp -3599
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp -3599
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp -3599
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp -3599
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp -3599
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp -3599
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_188
timestamp -3599
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_200
timestamp -3599
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636964856
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp -3599
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp -3599
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp -3599
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_237
timestamp -3599
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp -3599
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp -3599
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp -3599
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp -3599
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp -3599
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp -3599
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_287
timestamp -3599
transform 1 0 27508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_301
timestamp -3599
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp -3599
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_12
timestamp 1636964856
transform 1 0 2208 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_24
timestamp 1636964856
transform 1 0 3312 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_36
timestamp 1636964856
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp -3599
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636964856
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636964856
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636964856
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636964856
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp -3599
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -3599
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp -3599
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_121
timestamp -3599
transform 1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp -3599
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp -3599
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp -3599
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_209
timestamp -3599
transform 1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp -3599
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_228
timestamp -3599
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_232
timestamp -3599
transform 1 0 22448 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_264
timestamp 1636964856
transform 1 0 25392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp -3599
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636964856
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp -3599
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_299
timestamp -3599
transform 1 0 28612 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7
timestamp 1636964856
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp -3599
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -3599
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636964856
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636964856
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636964856
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636964856
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp -3599
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp -3599
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp -3599
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp -3599
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_98
timestamp -3599
transform 1 0 10120 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_127
timestamp -3599
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp -3599
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp -3599
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_171
timestamp -3599
transform 1 0 16836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp -3599
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp -3599
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp -3599
transform 1 0 20056 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp -3599
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636964856
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636964856
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636964856
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636964856
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_301
timestamp -3599
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636964856
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636964856
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636964856
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636964856
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp -3599
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp -3599
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636964856
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636964856
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_81
timestamp -3599
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_105
timestamp -3599
transform 1 0 10764 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp -3599
transform 1 0 12420 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_134
timestamp -3599
transform 1 0 13432 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp -3599
transform 1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_154
timestamp -3599
transform 1 0 15272 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_162
timestamp -3599
transform 1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_172
timestamp -3599
transform 1 0 16928 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_186
timestamp -3599
transform 1 0 18216 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_194
timestamp -3599
transform 1 0 18952 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_198
timestamp -3599
transform 1 0 19320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp -3599
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp -3599
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636964856
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_237
timestamp -3599
transform 1 0 22908 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1636964856
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp -3599
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp -3599
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636964856
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636964856
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_305
timestamp -3599
transform 1 0 29164 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636964856
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636964856
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -3599
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636964856
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636964856
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636964856
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636964856
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp -3599
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -3599
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636964856
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636964856
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp -3599
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_116
timestamp -3599
transform 1 0 11776 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_120
timestamp -3599
transform 1 0 12144 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_129
timestamp -3599
transform 1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp -3599
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_141
timestamp -3599
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_156
timestamp 1636964856
transform 1 0 15456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp -3599
transform 1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_173
timestamp 1636964856
transform 1 0 17020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp -3599
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636964856
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_212
timestamp 1636964856
transform 1 0 20608 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp -3599
transform 1 0 21712 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp -3599
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_253
timestamp -3599
transform 1 0 24380 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_257
timestamp 1636964856
transform 1 0 24748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_269
timestamp 1636964856
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1636964856
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1636964856
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp -3599
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1636964856
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1636964856
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_31
timestamp -3599
transform 1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp -3599
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -3599
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_80
timestamp -3599
transform 1 0 8464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_90
timestamp -3599
transform 1 0 9384 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_96
timestamp -3599
transform 1 0 9936 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_103
timestamp -3599
transform 1 0 10580 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_120
timestamp -3599
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp -3599
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp -3599
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp -3599
transform 1 0 16928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp -3599
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_202
timestamp -3599
transform 1 0 19688 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_212
timestamp -3599
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_222
timestamp -3599
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp -3599
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_236
timestamp -3599
transform 1 0 22816 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_244
timestamp -3599
transform 1 0 23552 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_250
timestamp 1636964856
transform 1 0 24104 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_262
timestamp 1636964856
transform 1 0 25208 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_274
timestamp -3599
transform 1 0 26312 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1636964856
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_293
timestamp -3599
transform 1 0 28060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_301
timestamp -3599
transform 1 0 28796 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636964856
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636964856
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -3599
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp -3599
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_54
timestamp -3599
transform 1 0 6072 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_69
timestamp -3599
transform 1 0 7452 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp -3599
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_96
timestamp -3599
transform 1 0 9936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp -3599
transform 1 0 11316 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_119
timestamp -3599
transform 1 0 12052 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_127
timestamp -3599
transform 1 0 12788 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp -3599
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp -3599
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_148
timestamp 1636964856
transform 1 0 14720 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_160
timestamp -3599
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_172
timestamp -3599
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp -3599
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp -3599
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_201
timestamp -3599
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp -3599
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp -3599
transform 1 0 21436 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_225
timestamp -3599
transform 1 0 21804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_238
timestamp 1636964856
transform 1 0 23000 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp -3599
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_260
timestamp 1636964856
transform 1 0 25024 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_272
timestamp 1636964856
transform 1 0 26128 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_284
timestamp 1636964856
transform 1 0 27232 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_296
timestamp 1636964856
transform 1 0 28336 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_16
timestamp 1636964856
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_28
timestamp 1636964856
transform 1 0 3680 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_40
timestamp 1636964856
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp -3599
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_64
timestamp 1636964856
transform 1 0 6992 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_83
timestamp 1636964856
transform 1 0 8740 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp -3599
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp -3599
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -3599
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_120
timestamp -3599
transform 1 0 12144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_126
timestamp -3599
transform 1 0 12696 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_132
timestamp -3599
transform 1 0 13248 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_142
timestamp -3599
transform 1 0 14168 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp -3599
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp -3599
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp -3599
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_178
timestamp 1636964856
transform 1 0 17480 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_190
timestamp 1636964856
transform 1 0 18584 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_202
timestamp -3599
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_213
timestamp -3599
transform 1 0 20700 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp -3599
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_232
timestamp -3599
transform 1 0 22448 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_264
timestamp 1636964856
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp -3599
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1636964856
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_293
timestamp -3599
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_297
timestamp -3599
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp -3599
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_29
timestamp -3599
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_33
timestamp -3599
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636964856
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636964856
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp -3599
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_79
timestamp -3599
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -3599
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_90
timestamp -3599
transform 1 0 9384 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_105
timestamp 1636964856
transform 1 0 10764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp -3599
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp -3599
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636964856
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_153
timestamp -3599
transform 1 0 15180 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_161
timestamp -3599
transform 1 0 15916 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp -3599
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_175
timestamp -3599
transform 1 0 17204 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp -3599
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_191
timestamp -3599
transform 1 0 18676 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp -3599
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1636964856
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_219
timestamp 1636964856
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_231
timestamp 1636964856
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_243
timestamp -3599
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp -3599
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1636964856
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1636964856
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1636964856
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1636964856
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp -3599
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp -3599
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636964856
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp -3599
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_42
timestamp -3599
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_46
timestamp -3599
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -3599
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_71
timestamp -3599
transform 1 0 7636 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_97
timestamp -3599
transform 1 0 10028 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp -3599
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_131
timestamp -3599
transform 1 0 13156 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp -3599
transform 1 0 13708 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_146
timestamp -3599
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_162
timestamp -3599
transform 1 0 16008 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_184
timestamp -3599
transform 1 0 18032 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_203
timestamp -3599
transform 1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp -3599
transform 1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp -3599
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp -3599
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636964856
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_256
timestamp 1636964856
transform 1 0 24656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_268
timestamp 1636964856
transform 1 0 25760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1636964856
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1636964856
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_305
timestamp -3599
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp -3599
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_17
timestamp -3599
transform 1 0 2668 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp -3599
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp -3599
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp -3599
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_46
timestamp -3599
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_57
timestamp -3599
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_66
timestamp -3599
transform 1 0 7176 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp -3599
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp -3599
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp -3599
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp -3599
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_99
timestamp -3599
transform 1 0 10212 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_114
timestamp -3599
transform 1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_122
timestamp -3599
transform 1 0 12328 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_131
timestamp -3599
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_150
timestamp -3599
transform 1 0 14904 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_159
timestamp 1636964856
transform 1 0 15732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp -3599
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_176
timestamp 1636964856
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp -3599
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp -3599
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_204
timestamp -3599
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_214
timestamp -3599
transform 1 0 20792 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_236
timestamp -3599
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_260
timestamp 1636964856
transform 1 0 25024 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_272
timestamp 1636964856
transform 1 0 26128 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_284
timestamp 1636964856
transform 1 0 27232 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_296
timestamp -3599
transform 1 0 28336 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_13
timestamp 1636964856
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_25
timestamp 1636964856
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_37
timestamp -3599
transform 1 0 4508 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp -3599
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_45
timestamp -3599
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp -3599
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp -3599
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_71
timestamp 1636964856
transform 1 0 7636 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_83
timestamp 1636964856
transform 1 0 8740 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_95
timestamp 1636964856
transform 1 0 9844 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp -3599
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -3599
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_116
timestamp -3599
transform 1 0 11776 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_128
timestamp -3599
transform 1 0 12880 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp -3599
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_141
timestamp -3599
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp -3599
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_175
timestamp -3599
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_179
timestamp 1636964856
transform 1 0 17572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_191
timestamp -3599
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_202
timestamp -3599
transform 1 0 19688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp -3599
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp -3599
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636964856
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp -3599
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_241
timestamp -3599
transform 1 0 23276 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_252
timestamp 1636964856
transform 1 0 24288 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_264
timestamp -3599
transform 1 0 25392 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_268
timestamp 1636964856
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1636964856
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_293
timestamp -3599
transform 1 0 28060 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_301
timestamp -3599
transform 1 0 28796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp -3599
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp -3599
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp -3599
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp -3599
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp -3599
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp -3599
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp -3599
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636964856
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_162
timestamp -3599
transform 1 0 16008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp -3599
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp -3599
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp -3599
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_220
timestamp -3599
transform 1 0 21344 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_237
timestamp -3599
transform 1 0 22908 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp -3599
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_253
timestamp -3599
transform 1 0 24380 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_257
timestamp 1636964856
transform 1 0 24748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_269
timestamp 1636964856
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_281
timestamp -3599
transform 1 0 26956 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_287
timestamp 1636964856
transform 1 0 27508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_299
timestamp -3599
transform 1 0 28612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp -3599
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_33
timestamp -3599
transform 1 0 4140 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp -3599
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp -3599
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp -3599
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_71
timestamp 1636964856
transform 1 0 7636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp -3599
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_99
timestamp 1636964856
transform 1 0 10212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -3599
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp -3599
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_126
timestamp -3599
transform 1 0 12696 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_134
timestamp -3599
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_139
timestamp -3599
transform 1 0 13892 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp -3599
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_152
timestamp 1636964856
transform 1 0 15088 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp -3599
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_179
timestamp 1636964856
transform 1 0 17572 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_191
timestamp 1636964856
transform 1 0 18676 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_203
timestamp 1636964856
transform 1 0 19780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_218
timestamp -3599
transform 1 0 21160 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp -3599
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_228
timestamp 1636964856
transform 1 0 22080 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_240
timestamp -3599
transform 1 0 23184 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_248
timestamp 1636964856
transform 1 0 23920 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_260
timestamp 1636964856
transform 1 0 25024 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp -3599
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_301
timestamp -3599
transform 1 0 28796 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636964856
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636964856
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -3599
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp -3599
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp -3599
transform 1 0 4692 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_44
timestamp 1636964856
transform 1 0 5152 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp -3599
transform 1 0 6256 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_67
timestamp -3599
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_76
timestamp -3599
transform 1 0 8096 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp -3599
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_107
timestamp -3599
transform 1 0 10948 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp -3599
transform 1 0 12880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_169
timestamp -3599
transform 1 0 16652 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_175
timestamp -3599
transform 1 0 17204 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_181
timestamp -3599
transform 1 0 17756 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp -3599
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp -3599
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_208
timestamp 1636964856
transform 1 0 20240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_220
timestamp -3599
transform 1 0 21344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_229
timestamp -3599
transform 1 0 22172 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp -3599
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_245
timestamp -3599
transform 1 0 23644 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636964856
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_265
timestamp -3599
transform 1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_275
timestamp -3599
transform 1 0 26404 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_283
timestamp -3599
transform 1 0 27140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_7
timestamp -3599
transform 1 0 1748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp -3599
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_32
timestamp -3599
transform 1 0 4048 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_40
timestamp -3599
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp -3599
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp -3599
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_57
timestamp -3599
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_66
timestamp -3599
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_93
timestamp -3599
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp -3599
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_143
timestamp 1636964856
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1636964856
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp -3599
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp -3599
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp -3599
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp -3599
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_185
timestamp -3599
transform 1 0 18124 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_191
timestamp -3599
transform 1 0 18676 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp -3599
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_205
timestamp -3599
transform 1 0 19964 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_211
timestamp -3599
transform 1 0 20516 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp -3599
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_228
timestamp -3599
transform 1 0 22080 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_259
timestamp -3599
transform 1 0 24932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp -3599
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_295
timestamp 1636964856
transform 1 0 28244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_307
timestamp -3599
transform 1 0 29348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp -3599
transform 1 0 2024 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_44
timestamp -3599
transform 1 0 5152 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_52
timestamp -3599
transform 1 0 5888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp -3599
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_95
timestamp -3599
transform 1 0 9844 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_105
timestamp -3599
transform 1 0 10764 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_120
timestamp -3599
transform 1 0 12144 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp -3599
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp -3599
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp -3599
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_170
timestamp -3599
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_182
timestamp -3599
transform 1 0 17848 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_190
timestamp -3599
transform 1 0 18584 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp -3599
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_242
timestamp -3599
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp -3599
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1636964856
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp -3599
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_275
timestamp -3599
transform 1 0 26404 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_283
timestamp -3599
transform 1 0 27140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_296
timestamp -3599
transform 1 0 28336 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_303
timestamp -3599
transform 1 0 28980 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636964856
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636964856
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636964856
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_39
timestamp -3599
transform 1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp -3599
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp -3599
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp -3599
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp -3599
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_79
timestamp -3599
transform 1 0 8372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp -3599
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp -3599
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_101
timestamp -3599
transform 1 0 10396 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp -3599
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp -3599
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_138
timestamp -3599
transform 1 0 13800 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_152
timestamp 1636964856
transform 1 0 15088 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp -3599
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp -3599
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_179
timestamp 1636964856
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp -3599
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_198
timestamp -3599
transform 1 0 19320 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp -3599
transform 1 0 20056 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp -3599
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp -3599
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_281
timestamp -3599
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp -3599
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp -3599
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp -3599
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_36
timestamp -3599
transform 1 0 4416 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_47
timestamp -3599
transform 1 0 5428 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_61
timestamp -3599
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_69
timestamp -3599
transform 1 0 7452 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp -3599
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp -3599
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp -3599
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_115
timestamp -3599
transform 1 0 11684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_123
timestamp -3599
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp -3599
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp -3599
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_153
timestamp -3599
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_157
timestamp -3599
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_161
timestamp 1636964856
transform 1 0 15916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp -3599
transform 1 0 17020 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_184
timestamp 1636964856
transform 1 0 18032 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_206
timestamp 1636964856
transform 1 0 20056 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_218
timestamp -3599
transform 1 0 21160 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp -3599
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_228
timestamp -3599
transform 1 0 22080 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp -3599
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_237
timestamp -3599
transform 1 0 22908 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp -3599
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp -3599
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_262
timestamp -3599
transform 1 0 25208 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_287
timestamp 1636964856
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp -3599
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp -3599
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_33
timestamp -3599
transform 1 0 4140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp -3599
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_64
timestamp -3599
transform 1 0 6992 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_76
timestamp -3599
transform 1 0 8096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_101
timestamp -3599
transform 1 0 10396 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_107
timestamp -3599
transform 1 0 10948 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -3599
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636964856
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636964856
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_137
timestamp -3599
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp -3599
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp -3599
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp -3599
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp -3599
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_228
timestamp 1636964856
transform 1 0 22080 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_240
timestamp 1636964856
transform 1 0 23184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_252
timestamp -3599
transform 1 0 24288 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_272
timestamp -3599
transform 1 0 26128 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_276
timestamp -3599
transform 1 0 26496 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp -3599
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_299
timestamp -3599
transform 1 0 28612 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_303
timestamp -3599
transform 1 0 28980 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp -3599
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp -3599
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_13
timestamp -3599
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_22
timestamp -3599
transform 1 0 3128 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_38
timestamp 1636964856
transform 1 0 4600 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_50
timestamp -3599
transform 1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_59
timestamp -3599
transform 1 0 6532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp -3599
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp -3599
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1636964856
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp -3599
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp -3599
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_109
timestamp -3599
transform 1 0 11132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_113
timestamp -3599
transform 1 0 11500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_125
timestamp -3599
transform 1 0 12604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_131
timestamp -3599
transform 1 0 13156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp -3599
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_141
timestamp -3599
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp -3599
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_174
timestamp -3599
transform 1 0 17112 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_183
timestamp 1636964856
transform 1 0 17940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp -3599
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636964856
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_233
timestamp -3599
transform 1 0 22540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_241
timestamp -3599
transform 1 0 23276 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp -3599
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_280
timestamp -3599
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_13
timestamp -3599
transform 1 0 2300 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp -3599
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp -3599
transform 1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp -3599
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -3599
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_65
timestamp -3599
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_72
timestamp 1636964856
transform 1 0 7728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_84
timestamp -3599
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_95
timestamp -3599
transform 1 0 9844 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -3599
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_126
timestamp -3599
transform 1 0 12696 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_148
timestamp -3599
transform 1 0 14720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp -3599
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp -3599
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_179
timestamp -3599
transform 1 0 17572 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_185
timestamp -3599
transform 1 0 18124 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_194
timestamp -3599
transform 1 0 18952 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp -3599
transform 1 0 19688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp -3599
transform 1 0 20608 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp -3599
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp -3599
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp -3599
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp -3599
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp -3599
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_289
timestamp 1636964856
transform 1 0 27692 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636964856
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp -3599
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp -3599
transform 1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_29
timestamp -3599
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp -3599
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_88
timestamp -3599
transform 1 0 9200 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_104
timestamp -3599
transform 1 0 10672 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1636964856
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_120
timestamp -3599
transform 1 0 12144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_128
timestamp -3599
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_135
timestamp -3599
transform 1 0 13524 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp -3599
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp -3599
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp -3599
transform 1 0 14812 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_155
timestamp -3599
transform 1 0 15364 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_166
timestamp 1636964856
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_188
timestamp -3599
transform 1 0 18400 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp -3599
transform 1 0 19504 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_225
timestamp 1636964856
transform 1 0 21804 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_237
timestamp 1636964856
transform 1 0 22908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_249
timestamp -3599
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp -3599
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp -3599
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_278
timestamp -3599
transform 1 0 26680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_282
timestamp -3599
transform 1 0 27048 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636964856
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636964856
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1636964856
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1636964856
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp -3599
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp -3599
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp -3599
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_66
timestamp 1636964856
transform 1 0 7176 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_78
timestamp 1636964856
transform 1 0 8280 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_90
timestamp -3599
transform 1 0 9384 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_99
timestamp 1636964856
transform 1 0 10212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp -3599
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_125
timestamp -3599
transform 1 0 12604 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_136
timestamp -3599
transform 1 0 13616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp -3599
transform 1 0 14168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp -3599
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp -3599
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_176
timestamp 1636964856
transform 1 0 17296 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_188
timestamp 1636964856
transform 1 0 18400 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_200
timestamp 1636964856
transform 1 0 19504 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_212
timestamp 1636964856
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_232
timestamp -3599
transform 1 0 22448 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_261
timestamp -3599
transform 1 0 25116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp -3599
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp -3599
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_300
timestamp -3599
transform 1 0 28704 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_7
timestamp -3599
transform 1 0 1748 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_18
timestamp -3599
transform 1 0 2760 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_24
timestamp -3599
transform 1 0 3312 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp -3599
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_38
timestamp -3599
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_50
timestamp -3599
transform 1 0 5704 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_58
timestamp -3599
transform 1 0 6440 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_68
timestamp 1636964856
transform 1 0 7360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp -3599
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_88
timestamp -3599
transform 1 0 9200 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_96
timestamp -3599
transform 1 0 9936 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_103
timestamp -3599
transform 1 0 10580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp -3599
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_117
timestamp -3599
transform 1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp -3599
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_175
timestamp -3599
transform 1 0 17204 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp -3599
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_206
timestamp -3599
transform 1 0 20056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_212
timestamp -3599
transform 1 0 20608 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_219
timestamp -3599
transform 1 0 21252 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_24_234
timestamp -3599
transform 1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_249
timestamp -3599
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_256
timestamp 1636964856
transform 1 0 24656 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_268
timestamp 1636964856
transform 1 0 25760 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_280
timestamp -3599
transform 1 0 26864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_284
timestamp -3599
transform 1 0 27232 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp -3599
transform 1 0 27600 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_296
timestamp -3599
transform 1 0 28336 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp -3599
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp -3599
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_49
timestamp -3599
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp -3599
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp -3599
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp -3599
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp -3599
transform 1 0 12420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_131
timestamp -3599
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp -3599
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp -3599
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_169
timestamp -3599
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_177
timestamp -3599
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_185
timestamp -3599
transform 1 0 18124 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_191
timestamp -3599
transform 1 0 18676 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_199
timestamp -3599
transform 1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp -3599
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_232
timestamp -3599
transform 1 0 22448 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp -3599
transform 1 0 24840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp -3599
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_271
timestamp -3599
transform 1 0 26036 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp -3599
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp -3599
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_7
timestamp 1636964856
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp -3599
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp -3599
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636964856
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1636964856
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_53
timestamp -3599
transform 1 0 5980 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_62
timestamp -3599
transform 1 0 6808 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp -3599
transform 1 0 7176 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_74
timestamp -3599
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp -3599
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636964856
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp -3599
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_102
timestamp -3599
transform 1 0 10488 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_108
timestamp 1636964856
transform 1 0 11040 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_120
timestamp -3599
transform 1 0 12144 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp -3599
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -3599
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp -3599
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_146
timestamp -3599
transform 1 0 14536 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp -3599
transform 1 0 15088 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_176
timestamp -3599
transform 1 0 17296 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp -3599
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp -3599
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636964856
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp -3599
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_227
timestamp -3599
transform 1 0 21988 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_237
timestamp 1636964856
transform 1 0 22908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp -3599
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp -3599
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_288
timestamp -3599
transform 1 0 27600 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_294
timestamp -3599
transform 1 0 28152 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_7
timestamp 1636964856
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_19
timestamp -3599
transform 1 0 2852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_28
timestamp -3599
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1636964856
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp -3599
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp -3599
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp -3599
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp -3599
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_74
timestamp -3599
transform 1 0 7912 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_90
timestamp -3599
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_96
timestamp -3599
transform 1 0 9936 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_108
timestamp -3599
transform 1 0 11040 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp -3599
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp -3599
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_133
timestamp -3599
transform 1 0 13340 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_147
timestamp 1636964856
transform 1 0 14628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp -3599
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_163
timestamp -3599
transform 1 0 16100 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp -3599
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636964856
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp -3599
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_191
timestamp -3599
transform 1 0 18676 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp -3599
transform 1 0 19780 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp -3599
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_213
timestamp -3599
transform 1 0 20700 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_233
timestamp 1636964856
transform 1 0 22540 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_245
timestamp 1636964856
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_257
timestamp -3599
transform 1 0 24748 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_263
timestamp -3599
transform 1 0 25300 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_269
timestamp -3599
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp -3599
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp -3599
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_306
timestamp -3599
transform 1 0 29256 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp -3599
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp -3599
transform 1 0 2116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_23
timestamp -3599
transform 1 0 3220 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -3599
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp -3599
transform 1 0 4416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_52
timestamp -3599
transform 1 0 5888 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp -3599
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_88
timestamp 1636964856
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_100
timestamp -3599
transform 1 0 10304 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_113
timestamp -3599
transform 1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_125
timestamp 1636964856
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp -3599
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1636964856
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_153
timestamp -3599
transform 1 0 15180 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp -3599
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_165
timestamp -3599
transform 1 0 16284 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_170
timestamp 1636964856
transform 1 0 16744 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_182
timestamp 1636964856
transform 1 0 17848 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp -3599
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_220
timestamp -3599
transform 1 0 21344 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_229
timestamp 1636964856
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp -3599
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp -3599
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_256
timestamp -3599
transform 1 0 24656 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_288
timestamp 1636964856
transform 1 0 27600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp -3599
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp -3599
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp -3599
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_8
timestamp -3599
transform 1 0 1840 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1636964856
transform 1 0 2576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_28
timestamp -3599
transform 1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_35
timestamp 1636964856
transform 1 0 4324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp -3599
transform 1 0 5428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp -3599
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1636964856
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1636964856
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1636964856
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_93
timestamp -3599
transform 1 0 9660 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_102
timestamp -3599
transform 1 0 10488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp -3599
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp -3599
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_140
timestamp -3599
transform 1 0 13984 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_148
timestamp -3599
transform 1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp -3599
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp -3599
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_192
timestamp 1636964856
transform 1 0 18768 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_204
timestamp -3599
transform 1 0 19872 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_212
timestamp -3599
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp -3599
transform 1 0 21160 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_232
timestamp -3599
transform 1 0 22448 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_268
timestamp -3599
transform 1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_272
timestamp -3599
transform 1 0 26128 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp -3599
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp -3599
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp -3599
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_16
timestamp 1636964856
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp -3599
transform 1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_70
timestamp -3599
transform 1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp -3599
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_88
timestamp -3599
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_103
timestamp 1636964856
transform 1 0 10580 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_115
timestamp 1636964856
transform 1 0 11684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_127
timestamp 1636964856
transform 1 0 12788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp -3599
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_155
timestamp -3599
transform 1 0 15364 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_161
timestamp -3599
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp -3599
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp -3599
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp -3599
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp -3599
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_210
timestamp -3599
transform 1 0 20424 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_221
timestamp -3599
transform 1 0 21436 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_237
timestamp 1636964856
transform 1 0 22908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp -3599
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636964856
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636964856
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp -3599
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_295
timestamp -3599
transform 1 0 28244 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_26
timestamp 1636964856
transform 1 0 3496 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_38
timestamp -3599
transform 1 0 4600 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_48
timestamp -3599
transform 1 0 5520 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp -3599
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_70
timestamp -3599
transform 1 0 7544 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp -3599
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_98
timestamp -3599
transform 1 0 10120 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_104
timestamp -3599
transform 1 0 10672 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp -3599
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp -3599
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_130
timestamp 1636964856
transform 1 0 13064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_142
timestamp -3599
transform 1 0 14168 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_152
timestamp 1636964856
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp -3599
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_176
timestamp -3599
transform 1 0 17296 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_187
timestamp -3599
transform 1 0 18308 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_195
timestamp -3599
transform 1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp -3599
transform 1 0 19872 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp -3599
transform 1 0 21068 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp -3599
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636964856
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_260
timestamp -3599
transform 1 0 25024 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_267
timestamp -3599
transform 1 0 25668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_272
timestamp -3599
transform 1 0 26128 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_291
timestamp -3599
transform 1 0 27876 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_299
timestamp -3599
transform 1 0 28612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp -3599
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_11
timestamp -3599
transform 1 0 2116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp -3599
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp -3599
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp -3599
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp -3599
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_39
timestamp 1636964856
transform 1 0 4692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_66
timestamp -3599
transform 1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp -3599
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_88
timestamp -3599
transform 1 0 9200 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp -3599
transform 1 0 10488 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_119
timestamp -3599
transform 1 0 12052 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp -3599
transform 1 0 12604 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp -3599
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp -3599
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 1636964856
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_173
timestamp -3599
transform 1 0 17020 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp -3599
transform 1 0 17572 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp -3599
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp -3599
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_213
timestamp -3599
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_230
timestamp 1636964856
transform 1 0 22264 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_242
timestamp -3599
transform 1 0 23368 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp -3599
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp -3599
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_286
timestamp -3599
transform 1 0 27416 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636964856
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp -3599
transform 1 0 2484 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_23
timestamp -3599
transform 1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_57
timestamp -3599
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_81
timestamp -3599
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_96
timestamp -3599
transform 1 0 9936 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp -3599
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp -3599
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_141
timestamp -3599
transform 1 0 14076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_156
timestamp -3599
transform 1 0 15456 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp -3599
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp -3599
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_209
timestamp -3599
transform 1 0 20332 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp -3599
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_225
timestamp -3599
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_231
timestamp -3599
transform 1 0 22356 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_258
timestamp 1636964856
transform 1 0 24840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_270
timestamp -3599
transform 1 0 25944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp -3599
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp -3599
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_292
timestamp 1636964856
transform 1 0 27968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_304
timestamp -3599
transform 1 0 29072 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1636964856
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1636964856
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp -3599
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp -3599
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_34
timestamp 1636964856
transform 1 0 4232 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_46
timestamp -3599
transform 1 0 5336 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp -3599
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp -3599
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_121
timestamp -3599
transform 1 0 12236 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp -3599
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp -3599
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636964856
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1636964856
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_165
timestamp -3599
transform 1 0 16284 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_174
timestamp -3599
transform 1 0 17112 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_180
timestamp -3599
transform 1 0 17664 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp -3599
transform 1 0 18308 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp -3599
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp -3599
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_241
timestamp -3599
transform 1 0 23276 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp -3599
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_287
timestamp 1636964856
transform 1 0 27508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_302
timestamp -3599
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1636964856
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_42
timestamp -3599
transform 1 0 4968 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp -3599
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_64
timestamp -3599
transform 1 0 6992 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_68
timestamp -3599
transform 1 0 7360 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_76
timestamp -3599
transform 1 0 8096 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp -3599
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_89
timestamp -3599
transform 1 0 9292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_93
timestamp -3599
transform 1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_101
timestamp -3599
transform 1 0 10396 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp -3599
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1636964856
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_125
timestamp -3599
transform 1 0 12604 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_134
timestamp -3599
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_142
timestamp -3599
transform 1 0 14168 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_158
timestamp -3599
transform 1 0 15640 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_179
timestamp -3599
transform 1 0 17572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_187
timestamp -3599
transform 1 0 18308 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_199
timestamp 1636964856
transform 1 0 19412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp -3599
transform 1 0 20516 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp -3599
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_228
timestamp -3599
transform 1 0 22080 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_236
timestamp -3599
transform 1 0 22816 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp -3599
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_307
timestamp -3599
transform 1 0 29348 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636964856
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636964856
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp -3599
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp -3599
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_39
timestamp 1636964856
transform 1 0 4692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp -3599
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_66
timestamp -3599
transform 1 0 7176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp -3599
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_101
timestamp -3599
transform 1 0 10396 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_127
timestamp -3599
transform 1 0 12788 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp -3599
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp -3599
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp -3599
transform 1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_156
timestamp 1636964856
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_168
timestamp -3599
transform 1 0 16560 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_174
timestamp 1636964856
transform 1 0 17112 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp -3599
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp -3599
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp -3599
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_209
timestamp -3599
transform 1 0 20332 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_238
timestamp -3599
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp -3599
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp -3599
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1636964856
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_299
timestamp -3599
transform 1 0 28612 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp -3599
transform 1 0 2300 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_17
timestamp -3599
transform 1 0 2668 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_44
timestamp -3599
transform 1 0 5152 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_60
timestamp -3599
transform 1 0 6624 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_75
timestamp -3599
transform 1 0 8004 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_83
timestamp -3599
transform 1 0 8740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_88
timestamp -3599
transform 1 0 9200 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_97
timestamp -3599
transform 1 0 10028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_104
timestamp -3599
transform 1 0 10672 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp -3599
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp -3599
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_117
timestamp -3599
transform 1 0 11868 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_132
timestamp 1636964856
transform 1 0 13248 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_144
timestamp 1636964856
transform 1 0 14352 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_156
timestamp 1636964856
transform 1 0 15456 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp -3599
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_201
timestamp -3599
transform 1 0 19596 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_219
timestamp -3599
transform 1 0 21252 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_265
timestamp 1636964856
transform 1 0 25484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_277
timestamp -3599
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_284
timestamp -3599
transform 1 0 27232 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636964856
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1636964856
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp -3599
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_29
timestamp -3599
transform 1 0 3772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_38
timestamp -3599
transform 1 0 4600 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1636964856
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_65
timestamp -3599
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_79
timestamp -3599
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp -3599
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1636964856
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp -3599
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_105
timestamp -3599
transform 1 0 10764 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_112
timestamp -3599
transform 1 0 11408 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_120
timestamp -3599
transform 1 0 12144 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_130
timestamp -3599
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp -3599
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_162
timestamp -3599
transform 1 0 16008 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp -3599
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636964856
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp -3599
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp -3599
transform 1 0 20700 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_241
timestamp -3599
transform 1 0 23276 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp -3599
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_262
timestamp 1636964856
transform 1 0 25208 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_274
timestamp -3599
transform 1 0 26312 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_282
timestamp -3599
transform 1 0 27048 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_296
timestamp 1636964856
transform 1 0 28336 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_13
timestamp -3599
transform 1 0 2300 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_21
timestamp -3599
transform 1 0 3036 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_25
timestamp -3599
transform 1 0 3404 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_43
timestamp -3599
transform 1 0 5060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_51
timestamp -3599
transform 1 0 5796 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp -3599
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_57
timestamp -3599
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_39_63
timestamp -3599
transform 1 0 6900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_74
timestamp -3599
transform 1 0 7912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_85
timestamp -3599
transform 1 0 8924 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_121
timestamp -3599
transform 1 0 12236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_136
timestamp -3599
transform 1 0 13616 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_146
timestamp 1636964856
transform 1 0 14536 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_158
timestamp -3599
transform 1 0 15640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp -3599
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_174
timestamp 1636964856
transform 1 0 17112 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_186
timestamp -3599
transform 1 0 18216 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_196
timestamp -3599
transform 1 0 19136 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_200
timestamp -3599
transform 1 0 19504 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_205
timestamp -3599
transform 1 0 19964 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_213
timestamp -3599
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_221
timestamp -3599
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636964856
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636964856
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636964856
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636964856
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_273
timestamp -3599
transform 1 0 26220 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_295
timestamp -3599
transform 1 0 28244 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp -3599
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_7
timestamp -3599
transform 1 0 1748 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp -3599
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_44
timestamp -3599
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_48
timestamp -3599
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_60
timestamp -3599
transform 1 0 6624 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_68
timestamp -3599
transform 1 0 7360 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_107
timestamp -3599
transform 1 0 10948 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_115
timestamp -3599
transform 1 0 11684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_132
timestamp -3599
transform 1 0 13248 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp -3599
transform 1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_161
timestamp -3599
transform 1 0 15916 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_179
timestamp -3599
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp -3599
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp -3599
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_230
timestamp -3599
transform 1 0 22264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_234
timestamp -3599
transform 1 0 22632 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_243
timestamp -3599
transform 1 0 23460 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp -3599
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_284
timestamp -3599
transform 1 0 27232 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_7
timestamp 1636964856
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_19
timestamp 1636964856
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1636964856
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_43
timestamp -3599
transform 1 0 5060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp -3599
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp -3599
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_66
timestamp -3599
transform 1 0 7176 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_77
timestamp 1636964856
transform 1 0 8188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_89
timestamp -3599
transform 1 0 9292 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_98
timestamp 1636964856
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp -3599
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1636964856
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1636964856
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp -3599
transform 1 0 13708 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_145
timestamp -3599
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_150
timestamp -3599
transform 1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_160
timestamp -3599
transform 1 0 15824 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_182
timestamp -3599
transform 1 0 17848 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_190
timestamp -3599
transform 1 0 18584 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_198
timestamp -3599
transform 1 0 19320 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_202
timestamp -3599
transform 1 0 19688 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_206
timestamp 1636964856
transform 1 0 20056 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp -3599
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_41_270
timestamp -3599
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp -3599
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_281
timestamp -3599
transform 1 0 26956 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_289
timestamp 1636964856
transform 1 0 27692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_301
timestamp -3599
transform 1 0 28796 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1636964856
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1636964856
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp -3599
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp -3599
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_40
timestamp 1636964856
transform 1 0 4784 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_52
timestamp -3599
transform 1 0 5888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_63
timestamp -3599
transform 1 0 6900 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_67
timestamp -3599
transform 1 0 7268 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_75
timestamp -3599
transform 1 0 8004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_79
timestamp -3599
transform 1 0 8372 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp -3599
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_85
timestamp -3599
transform 1 0 8924 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_89
timestamp -3599
transform 1 0 9292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp -3599
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_118
timestamp -3599
transform 1 0 11960 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp -3599
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp -3599
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_141
timestamp -3599
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_148
timestamp 1636964856
transform 1 0 14720 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_166
timestamp -3599
transform 1 0 16376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_170
timestamp -3599
transform 1 0 16744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_180
timestamp -3599
transform 1 0 17664 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp -3599
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp -3599
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp -3599
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_201
timestamp -3599
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_205
timestamp 1636964856
transform 1 0 19964 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_217
timestamp -3599
transform 1 0 21068 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_223
timestamp -3599
transform 1 0 21620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_232
timestamp -3599
transform 1 0 22448 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_246
timestamp -3599
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636964856
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636964856
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_277
timestamp -3599
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_283
timestamp -3599
transform 1 0 27140 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_287
timestamp -3599
transform 1 0 27508 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_293
timestamp -3599
transform 1 0 28060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_299
timestamp -3599
transform 1 0 28612 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_303
timestamp -3599
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp -3599
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636964856
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636964856
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_27
timestamp -3599
transform 1 0 3588 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_48
timestamp -3599
transform 1 0 5520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_57
timestamp -3599
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_67
timestamp -3599
transform 1 0 7268 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_81
timestamp -3599
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp -3599
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_124
timestamp -3599
transform 1 0 12512 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp -3599
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_160
timestamp -3599
transform 1 0 15824 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_175
timestamp -3599
transform 1 0 17204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_181
timestamp -3599
transform 1 0 17756 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_192
timestamp -3599
transform 1 0 18768 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_245
timestamp -3599
transform 1 0 23644 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_253
timestamp -3599
transform 1 0 24380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_259
timestamp -3599
transform 1 0 24932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp -3599
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp -3599
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_7
timestamp 1636964856
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp -3599
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp -3599
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_29
timestamp -3599
transform 1 0 3772 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_33
timestamp -3599
transform 1 0 4140 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_42
timestamp -3599
transform 1 0 4968 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_50
timestamp -3599
transform 1 0 5704 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_62
timestamp 1636964856
transform 1 0 6808 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_74
timestamp -3599
transform 1 0 7912 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp -3599
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp -3599
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_94
timestamp -3599
transform 1 0 9752 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_108
timestamp -3599
transform 1 0 11040 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_117
timestamp -3599
transform 1 0 11868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp -3599
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_141
timestamp -3599
transform 1 0 14076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_161
timestamp -3599
transform 1 0 15916 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_166
timestamp -3599
transform 1 0 16376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp -3599
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_200
timestamp -3599
transform 1 0 19504 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_214
timestamp 1636964856
transform 1 0 20792 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_226
timestamp 1636964856
transform 1 0 21896 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_238
timestamp -3599
transform 1 0 23000 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp -3599
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_293
timestamp -3599
transform 1 0 28060 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_301
timestamp -3599
transform 1 0 28796 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636964856
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636964856
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1636964856
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1636964856
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp -3599
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp -3599
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_62
timestamp -3599
transform 1 0 6808 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_66
timestamp -3599
transform 1 0 7176 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_72
timestamp -3599
transform 1 0 7728 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_97
timestamp 1636964856
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp -3599
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp -3599
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_121
timestamp -3599
transform 1 0 12236 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp -3599
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_131
timestamp -3599
transform 1 0 13156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_135
timestamp -3599
transform 1 0 13524 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_142
timestamp -3599
transform 1 0 14168 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_148
timestamp -3599
transform 1 0 14720 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_156
timestamp 1636964856
transform 1 0 15456 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1636964856
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_181
timestamp -3599
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_192
timestamp 1636964856
transform 1 0 18768 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_204
timestamp 1636964856
transform 1 0 19872 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_216
timestamp -3599
transform 1 0 20976 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp -3599
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp -3599
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_236
timestamp -3599
transform 1 0 22816 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_242
timestamp -3599
transform 1 0 23368 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_263
timestamp 1636964856
transform 1 0 25300 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_275
timestamp -3599
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp -3599
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp -3599
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_290
timestamp -3599
transform 1 0 27784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_298
timestamp -3599
transform 1 0 28520 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_13
timestamp 1636964856
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp -3599
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_29
timestamp -3599
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_37
timestamp -3599
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp -3599
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_88
timestamp -3599
transform 1 0 9200 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_94
timestamp -3599
transform 1 0 9752 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_98
timestamp -3599
transform 1 0 10120 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp -3599
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_141
timestamp -3599
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_153
timestamp -3599
transform 1 0 15180 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_161
timestamp -3599
transform 1 0 15916 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_169
timestamp -3599
transform 1 0 16652 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_175
timestamp -3599
transform 1 0 17204 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_185
timestamp -3599
transform 1 0 18124 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp -3599
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_253
timestamp -3599
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp -3599
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_271
timestamp 1636964856
transform 1 0 26036 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_283
timestamp -3599
transform 1 0 27140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp -3599
transform 1 0 27508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1636964856
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1636964856
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1636964856
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1636964856
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_54
timestamp -3599
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_60
timestamp 1636964856
transform 1 0 6624 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_103
timestamp -3599
transform 1 0 10580 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_110
timestamp -3599
transform 1 0 11224 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1636964856
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_153
timestamp -3599
transform 1 0 15180 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp -3599
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_190
timestamp -3599
transform 1 0 18584 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_206
timestamp -3599
transform 1 0 20056 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_214
timestamp -3599
transform 1 0 20792 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp -3599
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636964856
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_237
timestamp -3599
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_256
timestamp -3599
transform 1 0 24656 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_288
timestamp 1636964856
transform 1 0 27600 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_300
timestamp -3599
transform 1 0 28704 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636964856
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1636964856
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp -3599
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1636964856
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1636964856
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1636964856
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_65
timestamp -3599
transform 1 0 7084 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_78
timestamp -3599
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_48_88
timestamp -3599
transform 1 0 9200 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_96
timestamp -3599
transform 1 0 9936 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_121
timestamp -3599
transform 1 0 12236 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_131
timestamp -3599
transform 1 0 13156 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_135
timestamp -3599
transform 1 0 13524 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp -3599
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636964856
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_153
timestamp -3599
transform 1 0 15180 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_160
timestamp 1636964856
transform 1 0 15824 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_172
timestamp -3599
transform 1 0 16928 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_185
timestamp -3599
transform 1 0 18124 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_191
timestamp -3599
transform 1 0 18676 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp -3599
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_197
timestamp -3599
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_228
timestamp -3599
transform 1 0 22080 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636964856
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_269
timestamp 1636964856
transform 1 0 25852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_281
timestamp -3599
transform 1 0 26956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp -3599
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_23
timestamp 1636964856
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_35
timestamp 1636964856
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp -3599
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp -3599
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1636964856
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1636964856
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1636964856
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1636964856
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_105
timestamp -3599
transform 1 0 10764 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1636964856
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1636964856
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_137
timestamp -3599
transform 1 0 13708 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1636964856
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_202
timestamp 1636964856
transform 1 0 19688 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp -3599
transform 1 0 20792 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp -3599
transform 1 0 21528 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1636964856
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_237
timestamp -3599
transform 1 0 22908 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_242
timestamp 1636964856
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1636964856
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1636964856
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp -3599
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1636964856
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_293
timestamp -3599
transform 1 0 28060 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_301
timestamp -3599
transform 1 0 28796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_17
timestamp -3599
transform 1 0 2668 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp -3599
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1636964856
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1636964856
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1636964856
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1636964856
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp -3599
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp -3599
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1636964856
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1636964856
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1636964856
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1636964856
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp -3599
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1636964856
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1636964856
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1636964856
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1636964856
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp -3599
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp -3599
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1636964856
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1636964856
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1636964856
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1636964856
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp -3599
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp -3599
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1636964856
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1636964856
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1636964856
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_289
timestamp -3599
transform 1 0 27692 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_295
timestamp -3599
transform 1 0 28244 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_25
timestamp -3599
transform 1 0 3404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_29
timestamp -3599
transform 1 0 3772 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_34
timestamp -3599
transform 1 0 4232 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_42
timestamp -3599
transform 1 0 4968 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp -3599
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp -3599
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp -3599
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_65
timestamp -3599
transform 1 0 7084 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_69
timestamp -3599
transform 1 0 7452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_77
timestamp -3599
transform 1 0 8188 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_85
timestamp -3599
transform 1 0 8924 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_93
timestamp -3599
transform 1 0 9660 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_98
timestamp -3599
transform 1 0 10120 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_106
timestamp -3599
transform 1 0 10856 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp -3599
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_113
timestamp -3599
transform 1 0 11500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_121
timestamp -3599
transform 1 0 12236 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_125
timestamp -3599
transform 1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_133
timestamp -3599
transform 1 0 13340 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_139
timestamp -3599
transform 1 0 13892 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_141
timestamp -3599
transform 1 0 14076 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_149
timestamp -3599
transform 1 0 14812 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_153
timestamp -3599
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp -3599
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp -3599
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_169
timestamp -3599
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_181
timestamp -3599
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_188
timestamp -3599
transform 1 0 18400 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_197
timestamp -3599
transform 1 0 19228 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_203
timestamp -3599
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_211
timestamp -3599
transform 1 0 20516 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp -3599
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp -3599
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp -3599
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_231
timestamp -3599
transform 1 0 22356 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_237
timestamp -3599
transform 1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_245
timestamp -3599
transform 1 0 23644 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_253
timestamp -3599
transform 1 0 24380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_261
timestamp -3599
transform 1 0 25116 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_266
timestamp 1636964856
transform 1 0 25576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp -3599
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp -3599
transform 1 0 8464 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp -3599
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp -3599
transform -1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp -3599
transform -1 0 15916 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp -3599
transform 1 0 1380 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp -3599
transform -1 0 29440 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3599
transform 1 0 1748 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp -3599
transform -1 0 19780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp -3599
transform 1 0 1380 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp -3599
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp -3599
transform -1 0 29440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp -3599
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp -3599
transform 1 0 1380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input14
timestamp -3599
transform -1 0 29440 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -3599
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp -3599
transform -1 0 29440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp -3599
transform 1 0 1380 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp -3599
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp -3599
transform 1 0 26956 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp -3599
transform -1 0 28796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp -3599
transform -1 0 29440 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp -3599
transform -1 0 29440 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp -3599
transform -1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp -3599
transform 1 0 2668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp -3599
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp -3599
transform 1 0 21988 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp -3599
transform 1 0 12972 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp -3599
transform -1 0 29440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp -3599
transform -1 0 28704 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp -3599
transform 1 0 7176 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp -3599
transform 1 0 3772 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp -3599
transform 1 0 1380 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp -3599
transform -1 0 29440 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp -3599
transform -1 0 25576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp -3599
transform -1 0 29440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input36
timestamp -3599
transform -1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp -3599
transform -1 0 29440 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input38
timestamp -3599
transform -1 0 29440 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp -3599
transform 1 0 9752 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input40
timestamp -3599
transform 1 0 11040 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp -3599
transform -1 0 29440 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp -3599
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input43
timestamp -3599
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp -3599
transform -1 0 29440 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp -3599
transform -1 0 29440 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp -3599
transform 1 0 16836 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp -3599
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input48
timestamp -3599
transform 1 0 7176 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp -3599
transform -1 0 12604 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp -3599
transform -1 0 29440 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp -3599
transform -1 0 29072 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input52
timestamp -3599
transform 1 0 14904 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input53
timestamp -3599
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp -3599
transform -1 0 29440 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp -3599
transform -1 0 29440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp -3599
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input57
timestamp -3599
transform 1 0 18124 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp -3599
transform 1 0 5244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp -3599
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp -3599
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input61
timestamp -3599
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp -3599
transform 1 0 2024 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input63
timestamp -3599
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp -3599
transform -1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input65
timestamp -3599
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp -3599
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp -3599
transform -1 0 29440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp -3599
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp -3599
transform -1 0 29440 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp -3599
transform -1 0 29440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp -3599
transform -1 0 26220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp -3599
transform -1 0 29440 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp -3599
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp -3599
transform 1 0 1380 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp -3599
transform 1 0 1380 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp -3599
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp -3599
transform -1 0 19136 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input78
timestamp -3599
transform 1 0 3956 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp -3599
transform 1 0 13616 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp -3599
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp -3599
transform 1 0 2300 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp -3599
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input83
timestamp -3599
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp -3599
transform -1 0 28244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp -3599
transform -1 0 21068 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp -3599
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input87
timestamp -3599
transform -1 0 28520 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp -3599
transform -1 0 29440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp -3599
transform 1 0 3036 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp -3599
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input91
timestamp -3599
transform -1 0 6256 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input92
timestamp -3599
transform 1 0 10396 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input93
timestamp -3599
transform -1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp -3599
transform -1 0 29440 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp -3599
transform 1 0 17480 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input96
timestamp -3599
transform 1 0 23920 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input97
timestamp -3599
transform 1 0 22632 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp -3599
transform 1 0 2300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input99
timestamp -3599
transform 1 0 1380 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  output100
timestamp -3599
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output101
timestamp -3599
transform 1 0 29164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output102
timestamp -3599
transform 1 0 28244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_52
timestamp -3599
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3599
transform -1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_53
timestamp -3599
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3599
transform -1 0 29716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_54
timestamp -3599
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3599
transform -1 0 29716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_55
timestamp -3599
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3599
transform -1 0 29716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_56
timestamp -3599
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3599
transform -1 0 29716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_57
timestamp -3599
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3599
transform -1 0 29716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_58
timestamp -3599
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3599
transform -1 0 29716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_59
timestamp -3599
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3599
transform -1 0 29716 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_60
timestamp -3599
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3599
transform -1 0 29716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_61
timestamp -3599
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3599
transform -1 0 29716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_62
timestamp -3599
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3599
transform -1 0 29716 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_63
timestamp -3599
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3599
transform -1 0 29716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_64
timestamp -3599
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3599
transform -1 0 29716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_65
timestamp -3599
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3599
transform -1 0 29716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_66
timestamp -3599
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3599
transform -1 0 29716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_67
timestamp -3599
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3599
transform -1 0 29716 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_68
timestamp -3599
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3599
transform -1 0 29716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_69
timestamp -3599
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3599
transform -1 0 29716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_70
timestamp -3599
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3599
transform -1 0 29716 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_71
timestamp -3599
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3599
transform -1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_72
timestamp -3599
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3599
transform -1 0 29716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_73
timestamp -3599
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3599
transform -1 0 29716 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_74
timestamp -3599
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3599
transform -1 0 29716 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_75
timestamp -3599
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3599
transform -1 0 29716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_76
timestamp -3599
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3599
transform -1 0 29716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_77
timestamp -3599
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3599
transform -1 0 29716 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_78
timestamp -3599
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3599
transform -1 0 29716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_79
timestamp -3599
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3599
transform -1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_80
timestamp -3599
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3599
transform -1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_81
timestamp -3599
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3599
transform -1 0 29716 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_82
timestamp -3599
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3599
transform -1 0 29716 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_83
timestamp -3599
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3599
transform -1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_84
timestamp -3599
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3599
transform -1 0 29716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_85
timestamp -3599
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3599
transform -1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_86
timestamp -3599
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp -3599
transform -1 0 29716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_87
timestamp -3599
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp -3599
transform -1 0 29716 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_88
timestamp -3599
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp -3599
transform -1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_89
timestamp -3599
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp -3599
transform -1 0 29716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_90
timestamp -3599
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp -3599
transform -1 0 29716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_91
timestamp -3599
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp -3599
transform -1 0 29716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_92
timestamp -3599
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp -3599
transform -1 0 29716 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_93
timestamp -3599
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp -3599
transform -1 0 29716 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_94
timestamp -3599
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp -3599
transform -1 0 29716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_95
timestamp -3599
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp -3599
transform -1 0 29716 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_96
timestamp -3599
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp -3599
transform -1 0 29716 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_97
timestamp -3599
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp -3599
transform -1 0 29716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_98
timestamp -3599
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp -3599
transform -1 0 29716 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_99
timestamp -3599
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp -3599
transform -1 0 29716 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_100
timestamp -3599
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp -3599
transform -1 0 29716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_101
timestamp -3599
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp -3599
transform -1 0 29716 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_102
timestamp -3599
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp -3599
transform -1 0 29716 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_103
timestamp -3599
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp -3599
transform -1 0 29716 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp -3599
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp -3599
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp -3599
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp -3599
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_108
timestamp -3599
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_109
timestamp -3599
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_110
timestamp -3599
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_111
timestamp -3599
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_112
timestamp -3599
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_113
timestamp -3599
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_114
timestamp -3599
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_115
timestamp -3599
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_116
timestamp -3599
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_117
timestamp -3599
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_118
timestamp -3599
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_119
timestamp -3599
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_120
timestamp -3599
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_121
timestamp -3599
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_122
timestamp -3599
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_123
timestamp -3599
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_124
timestamp -3599
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_125
timestamp -3599
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_126
timestamp -3599
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_127
timestamp -3599
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_128
timestamp -3599
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_129
timestamp -3599
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_130
timestamp -3599
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_131
timestamp -3599
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_132
timestamp -3599
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_133
timestamp -3599
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_134
timestamp -3599
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_135
timestamp -3599
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_136
timestamp -3599
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_137
timestamp -3599
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_138
timestamp -3599
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_139
timestamp -3599
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_140
timestamp -3599
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_141
timestamp -3599
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_142
timestamp -3599
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_143
timestamp -3599
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_144
timestamp -3599
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_145
timestamp -3599
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_146
timestamp -3599
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_147
timestamp -3599
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_148
timestamp -3599
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_149
timestamp -3599
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_150
timestamp -3599
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_151
timestamp -3599
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_152
timestamp -3599
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_153
timestamp -3599
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_154
timestamp -3599
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_155
timestamp -3599
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_156
timestamp -3599
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_157
timestamp -3599
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_158
timestamp -3599
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_159
timestamp -3599
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_160
timestamp -3599
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_161
timestamp -3599
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_162
timestamp -3599
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_163
timestamp -3599
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_164
timestamp -3599
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_165
timestamp -3599
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_166
timestamp -3599
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_167
timestamp -3599
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_168
timestamp -3599
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_169
timestamp -3599
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_170
timestamp -3599
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_171
timestamp -3599
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_172
timestamp -3599
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_173
timestamp -3599
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_174
timestamp -3599
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_175
timestamp -3599
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_176
timestamp -3599
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_177
timestamp -3599
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_178
timestamp -3599
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_179
timestamp -3599
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_180
timestamp -3599
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_181
timestamp -3599
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_182
timestamp -3599
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_183
timestamp -3599
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_184
timestamp -3599
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_185
timestamp -3599
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_186
timestamp -3599
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_187
timestamp -3599
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_188
timestamp -3599
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_189
timestamp -3599
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_190
timestamp -3599
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_191
timestamp -3599
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_192
timestamp -3599
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_193
timestamp -3599
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_194
timestamp -3599
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_195
timestamp -3599
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_196
timestamp -3599
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_197
timestamp -3599
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_198
timestamp -3599
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_199
timestamp -3599
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_200
timestamp -3599
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_201
timestamp -3599
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_202
timestamp -3599
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_203
timestamp -3599
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_204
timestamp -3599
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_205
timestamp -3599
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_206
timestamp -3599
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_207
timestamp -3599
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_208
timestamp -3599
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_209
timestamp -3599
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_210
timestamp -3599
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_211
timestamp -3599
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_212
timestamp -3599
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_213
timestamp -3599
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_214
timestamp -3599
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_215
timestamp -3599
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_216
timestamp -3599
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_217
timestamp -3599
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_218
timestamp -3599
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_219
timestamp -3599
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_220
timestamp -3599
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_221
timestamp -3599
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_222
timestamp -3599
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_223
timestamp -3599
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_224
timestamp -3599
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_225
timestamp -3599
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_226
timestamp -3599
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_227
timestamp -3599
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_228
timestamp -3599
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_229
timestamp -3599
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_230
timestamp -3599
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_231
timestamp -3599
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_232
timestamp -3599
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_233
timestamp -3599
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_234
timestamp -3599
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_235
timestamp -3599
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_236
timestamp -3599
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_237
timestamp -3599
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_238
timestamp -3599
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_239
timestamp -3599
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_240
timestamp -3599
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_241
timestamp -3599
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_242
timestamp -3599
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_243
timestamp -3599
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_244
timestamp -3599
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_245
timestamp -3599
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_246
timestamp -3599
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_247
timestamp -3599
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_248
timestamp -3599
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_249
timestamp -3599
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_250
timestamp -3599
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_251
timestamp -3599
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_252
timestamp -3599
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_253
timestamp -3599
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_254
timestamp -3599
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_255
timestamp -3599
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_256
timestamp -3599
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_257
timestamp -3599
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_258
timestamp -3599
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_259
timestamp -3599
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_260
timestamp -3599
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_261
timestamp -3599
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_262
timestamp -3599
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_263
timestamp -3599
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_264
timestamp -3599
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_265
timestamp -3599
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_266
timestamp -3599
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_267
timestamp -3599
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_268
timestamp -3599
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_269
timestamp -3599
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_270
timestamp -3599
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_271
timestamp -3599
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_272
timestamp -3599
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_273
timestamp -3599
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_274
timestamp -3599
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_275
timestamp -3599
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_276
timestamp -3599
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_277
timestamp -3599
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_278
timestamp -3599
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_279
timestamp -3599
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_280
timestamp -3599
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_281
timestamp -3599
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_282
timestamp -3599
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_283
timestamp -3599
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_284
timestamp -3599
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_285
timestamp -3599
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_286
timestamp -3599
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_287
timestamp -3599
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_288
timestamp -3599
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_289
timestamp -3599
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_290
timestamp -3599
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_291
timestamp -3599
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_292
timestamp -3599
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_293
timestamp -3599
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_294
timestamp -3599
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_295
timestamp -3599
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_296
timestamp -3599
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_297
timestamp -3599
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_298
timestamp -3599
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp -3599
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp -3599
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp -3599
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp -3599
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_303
timestamp -3599
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_304
timestamp -3599
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_305
timestamp -3599
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_306
timestamp -3599
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_307
timestamp -3599
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_308
timestamp -3599
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_309
timestamp -3599
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_310
timestamp -3599
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_311
timestamp -3599
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_312
timestamp -3599
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_313
timestamp -3599
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_314
timestamp -3599
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_315
timestamp -3599
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_316
timestamp -3599
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_317
timestamp -3599
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_318
timestamp -3599
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_319
timestamp -3599
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_320
timestamp -3599
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_321
timestamp -3599
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_322
timestamp -3599
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_323
timestamp -3599
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_324
timestamp -3599
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_325
timestamp -3599
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_326
timestamp -3599
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_327
timestamp -3599
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_328
timestamp -3599
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_329
timestamp -3599
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_330
timestamp -3599
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_331
timestamp -3599
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_332
timestamp -3599
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_333
timestamp -3599
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_334
timestamp -3599
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_335
timestamp -3599
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_336
timestamp -3599
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_337
timestamp -3599
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_338
timestamp -3599
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_339
timestamp -3599
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_340
timestamp -3599
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_341
timestamp -3599
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_342
timestamp -3599
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_343
timestamp -3599
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_344
timestamp -3599
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_345
timestamp -3599
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_346
timestamp -3599
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_347
timestamp -3599
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_348
timestamp -3599
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp -3599
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_350
timestamp -3599
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_351
timestamp -3599
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_352
timestamp -3599
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_353
timestamp -3599
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_354
timestamp -3599
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_355
timestamp -3599
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_356
timestamp -3599
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_357
timestamp -3599
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_358
timestamp -3599
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_359
timestamp -3599
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_360
timestamp -3599
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_361
timestamp -3599
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_362
timestamp -3599
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_363
timestamp -3599
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_364
timestamp -3599
transform 1 0 3680 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_365
timestamp -3599
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_366
timestamp -3599
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_367
timestamp -3599
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_368
timestamp -3599
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_369
timestamp -3599
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_370
timestamp -3599
transform 1 0 19136 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_371
timestamp -3599
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_372
timestamp -3599
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_373
timestamp -3599
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
<< labels >>
flabel metal2 s 8390 32247 8446 33047 0 FreeSans 224 90 0 0 PWM_CNTA[0]
port 0 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 PWM_CNTA[10]
port 1 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 PWM_CNTA[11]
port 2 nsew signal input
flabel metal2 s 15474 32247 15530 33047 0 FreeSans 224 90 0 0 PWM_CNTA[12]
port 3 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 PWM_CNTA[13]
port 4 nsew signal input
flabel metal3 s 30103 12248 30903 12368 0 FreeSans 480 0 0 0 PWM_CNTA[14]
port 5 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 PWM_CNTA[15]
port 6 nsew signal input
flabel metal2 s 19338 32247 19394 33047 0 FreeSans 224 90 0 0 PWM_CNTA[16]
port 7 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 PWM_CNTA[17]
port 8 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 PWM_CNTA[18]
port 9 nsew signal input
flabel metal3 s 30103 25848 30903 25968 0 FreeSans 480 0 0 0 PWM_CNTA[19]
port 10 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 PWM_CNTA[1]
port 11 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 PWM_CNTA[20]
port 12 nsew signal input
flabel metal3 s 30103 7488 30903 7608 0 FreeSans 480 0 0 0 PWM_CNTA[21]
port 13 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 PWM_CNTA[22]
port 14 nsew signal input
flabel metal3 s 30103 17008 30903 17128 0 FreeSans 480 0 0 0 PWM_CNTA[23]
port 15 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 PWM_CNTA[24]
port 16 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 PWM_CNTA[25]
port 17 nsew signal input
flabel metal2 s 26422 32247 26478 33047 0 FreeSans 224 90 0 0 PWM_CNTA[26]
port 18 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 PWM_CNTA[27]
port 19 nsew signal input
flabel metal3 s 30103 6128 30903 6248 0 FreeSans 480 0 0 0 PWM_CNTA[28]
port 20 nsew signal input
flabel metal3 s 30103 18368 30903 18488 0 FreeSans 480 0 0 0 PWM_CNTA[29]
port 21 nsew signal input
flabel metal3 s 30103 29928 30903 30048 0 FreeSans 480 0 0 0 PWM_CNTA[2]
port 22 nsew signal input
flabel metal2 s 2594 32247 2650 33047 0 FreeSans 224 90 0 0 PWM_CNTA[30]
port 23 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 PWM_CNTA[31]
port 24 nsew signal input
flabel metal2 s 21914 32247 21970 33047 0 FreeSans 224 90 0 0 PWM_CNTA[3]
port 25 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 PWM_CNTA[4]
port 26 nsew signal input
flabel metal2 s 28998 32247 29054 33047 0 FreeSans 224 90 0 0 PWM_CNTA[5]
port 27 nsew signal input
flabel metal3 s 30103 31288 30903 31408 0 FreeSans 480 0 0 0 PWM_CNTA[6]
port 28 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 PWM_CNTA[7]
port 29 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 PWM_CNTA[8]
port 30 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 PWM_CNTA[9]
port 31 nsew signal input
flabel metal3 s 30103 32648 30903 32768 0 FreeSans 480 0 0 0 PWM_CNTB[0]
port 32 nsew signal input
flabel metal2 s 25134 32247 25190 33047 0 FreeSans 224 90 0 0 PWM_CNTB[10]
port 33 nsew signal input
flabel metal3 s 30103 2048 30903 2168 0 FreeSans 480 0 0 0 PWM_CNTB[11]
port 34 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 PWM_CNTB[12]
port 35 nsew signal input
flabel metal3 s 30103 14968 30903 15088 0 FreeSans 480 0 0 0 PWM_CNTB[13]
port 36 nsew signal input
flabel metal3 s 30103 10888 30903 11008 0 FreeSans 480 0 0 0 PWM_CNTB[14]
port 37 nsew signal input
flabel metal2 s 9678 32247 9734 33047 0 FreeSans 224 90 0 0 PWM_CNTB[15]
port 38 nsew signal input
flabel metal2 s 10966 32247 11022 33047 0 FreeSans 224 90 0 0 PWM_CNTB[16]
port 39 nsew signal input
flabel metal3 s 30103 24488 30903 24608 0 FreeSans 480 0 0 0 PWM_CNTB[17]
port 40 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 PWM_CNTB[18]
port 41 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 PWM_CNTB[19]
port 42 nsew signal input
flabel metal3 s 30103 27208 30903 27328 0 FreeSans 480 0 0 0 PWM_CNTB[1]
port 43 nsew signal input
flabel metal3 s 30103 688 30903 808 0 FreeSans 480 0 0 0 PWM_CNTB[20]
port 44 nsew signal input
flabel metal2 s 16762 32247 16818 33047 0 FreeSans 224 90 0 0 PWM_CNTB[21]
port 45 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 PWM_CNTB[22]
port 46 nsew signal input
flabel metal2 s 7102 32247 7158 33047 0 FreeSans 224 90 0 0 PWM_CNTB[23]
port 47 nsew signal input
flabel metal2 s 12254 32247 12310 33047 0 FreeSans 224 90 0 0 PWM_CNTB[24]
port 48 nsew signal input
flabel metal3 s 30103 28568 30903 28688 0 FreeSans 480 0 0 0 PWM_CNTB[25]
port 49 nsew signal input
flabel metal3 s 30103 8 30903 128 0 FreeSans 480 0 0 0 PWM_CNTB[26]
port 50 nsew signal input
flabel metal2 s 14830 32247 14886 33047 0 FreeSans 224 90 0 0 PWM_CNTB[27]
port 51 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 PWM_CNTB[28]
port 52 nsew signal input
flabel metal3 s 30103 8168 30903 8288 0 FreeSans 480 0 0 0 PWM_CNTB[29]
port 53 nsew signal input
flabel metal3 s 30103 21088 30903 21208 0 FreeSans 480 0 0 0 PWM_CNTB[2]
port 54 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 PWM_CNTB[30]
port 55 nsew signal input
flabel metal2 s 18050 32247 18106 33047 0 FreeSans 224 90 0 0 PWM_CNTB[31]
port 56 nsew signal input
flabel metal2 s 5170 32247 5226 33047 0 FreeSans 224 90 0 0 PWM_CNTB[3]
port 57 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 PWM_CNTB[4]
port 58 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 PWM_CNTB[5]
port 59 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 PWM_CNTB[6]
port 60 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 PWM_CNTB[7]
port 61 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 PWM_CNTB[8]
port 62 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 PWM_CNTB[9]
port 63 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 PWM_OUTA
port 64 nsew signal output
flabel metal3 s 30103 9528 30903 9648 0 FreeSans 480 0 0 0 PWM_OUTB
port 65 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 TIMER_TOP[0]
port 66 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 TIMER_TOP[10]
port 67 nsew signal input
flabel metal3 s 30103 3408 30903 3528 0 FreeSans 480 0 0 0 TIMER_TOP[11]
port 68 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 TIMER_TOP[12]
port 69 nsew signal input
flabel metal3 s 30103 13608 30903 13728 0 FreeSans 480 0 0 0 TIMER_TOP[13]
port 70 nsew signal input
flabel metal3 s 30103 22448 30903 22568 0 FreeSans 480 0 0 0 TIMER_TOP[14]
port 71 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 TIMER_TOP[15]
port 72 nsew signal input
flabel metal3 s 30103 23808 30903 23928 0 FreeSans 480 0 0 0 TIMER_TOP[16]
port 73 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 TIMER_TOP[17]
port 74 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 TIMER_TOP[18]
port 75 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 TIMER_TOP[19]
port 76 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 TIMER_TOP[1]
port 77 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 TIMER_TOP[20]
port 78 nsew signal input
flabel metal2 s 3882 32247 3938 33047 0 FreeSans 224 90 0 0 TIMER_TOP[21]
port 79 nsew signal input
flabel metal2 s 13542 32247 13598 33047 0 FreeSans 224 90 0 0 TIMER_TOP[22]
port 80 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 TIMER_TOP[23]
port 81 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 TIMER_TOP[24]
port 82 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 TIMER_TOP[25]
port 83 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 TIMER_TOP[26]
port 84 nsew signal input
flabel metal2 s 27710 32247 27766 33047 0 FreeSans 224 90 0 0 TIMER_TOP[27]
port 85 nsew signal input
flabel metal2 s 20626 32247 20682 33047 0 FreeSans 224 90 0 0 TIMER_TOP[28]
port 86 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 TIMER_TOP[29]
port 87 nsew signal input
flabel metal2 s 30286 32247 30342 33047 0 FreeSans 224 90 0 0 TIMER_TOP[2]
port 88 nsew signal input
flabel metal3 s 30103 4768 30903 4888 0 FreeSans 480 0 0 0 TIMER_TOP[30]
port 89 nsew signal input
flabel metal2 s 18 32247 74 33047 0 FreeSans 224 90 0 0 TIMER_TOP[31]
port 90 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 TIMER_TOP[3]
port 91 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 TIMER_TOP[4]
port 92 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 TIMER_TOP[5]
port 93 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 TIMER_TOP[6]
port 94 nsew signal input
flabel metal3 s 30103 19728 30903 19848 0 FreeSans 480 0 0 0 TIMER_TOP[7]
port 95 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 TIMER_TOP[8]
port 96 nsew signal input
flabel metal2 s 23846 32247 23902 33047 0 FreeSans 224 90 0 0 TIMER_TOP[9]
port 97 nsew signal input
flabel metal2 s 22558 32247 22614 33047 0 FreeSans 224 90 0 0 TMR_MODE[0]
port 98 nsew signal input
flabel metal2 s 1306 32247 1362 33047 0 FreeSans 224 90 0 0 TMR_MODE[1]
port 99 nsew signal input
flabel metal2 s 6458 32247 6514 33047 0 FreeSans 224 90 0 0 TMR_SRC[0]
port 100 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 TMR_SRC[1]
port 101 nsew signal input
flabel metal4 s 4868 2128 5188 30512 0 FreeSans 1920 90 0 0 VGND
port 102 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 30512 0 FreeSans 1920 90 0 0 VPWR
port 103 nsew power bidirectional
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 clk
port 104 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 reset
port 105 nsew signal input
flabel metal3 s 30103 16328 30903 16448 0 FreeSans 480 0 0 0 timer_interrupt
port 106 nsew signal output
rlabel metal1 15410 30464 15410 30464 0 VGND
rlabel metal1 15410 29920 15410 29920 0 VPWR
rlabel metal1 8510 30294 8510 30294 0 PWM_CNTA[0]
rlabel metal3 751 21148 751 21148 0 PWM_CNTA[10]
rlabel metal2 27094 1554 27094 1554 0 PWM_CNTA[11]
rlabel metal1 15640 30294 15640 30294 0 PWM_CNTA[12]
rlabel metal3 751 29988 751 29988 0 PWM_CNTA[13]
rlabel metal3 29770 12308 29770 12308 0 PWM_CNTA[14]
rlabel metal3 820 2108 820 2108 0 PWM_CNTA[15]
rlabel metal1 19504 30294 19504 30294 0 PWM_CNTA[16]
rlabel metal3 751 22508 751 22508 0 PWM_CNTA[17]
rlabel metal3 751 10948 751 10948 0 PWM_CNTA[18]
rlabel metal2 29302 26095 29302 26095 0 PWM_CNTA[19]
rlabel metal3 751 24548 751 24548 0 PWM_CNTA[1]
rlabel metal3 751 18428 751 18428 0 PWM_CNTA[20]
rlabel metal2 29394 7701 29394 7701 0 PWM_CNTA[21]
rlabel metal3 1096 15028 1096 15028 0 PWM_CNTA[22]
rlabel metal2 29302 16813 29302 16813 0 PWM_CNTA[23]
rlabel metal3 751 27268 751 27268 0 PWM_CNTA[24]
rlabel metal3 751 17068 751 17068 0 PWM_CNTA[25]
rlabel metal1 26726 30226 26726 30226 0 PWM_CNTA[26]
rlabel metal2 28382 1554 28382 1554 0 PWM_CNTA[27]
rlabel via2 29394 6205 29394 6205 0 PWM_CNTA[28]
rlabel metal2 29394 18581 29394 18581 0 PWM_CNTA[29]
rlabel metal2 28934 29801 28934 29801 0 PWM_CNTA[2]
rlabel metal2 2622 31290 2622 31290 0 PWM_CNTA[30]
rlabel metal3 751 19788 751 19788 0 PWM_CNTA[31]
rlabel metal2 21942 31290 21942 31290 0 PWM_CNTA[3]
rlabel metal2 12926 1588 12926 1588 0 PWM_CNTA[4]
rlabel metal1 29164 29614 29164 29614 0 PWM_CNTA[5]
rlabel metal2 28566 30481 28566 30481 0 PWM_CNTA[6]
rlabel metal2 7130 1588 7130 1588 0 PWM_CNTA[7]
rlabel metal2 3266 1588 3266 1588 0 PWM_CNTA[8]
rlabel metal3 751 6188 751 6188 0 PWM_CNTA[9]
rlabel metal2 29394 31467 29394 31467 0 PWM_CNTB[0]
rlabel metal1 25300 30294 25300 30294 0 PWM_CNTB[10]
rlabel metal2 29302 2227 29302 2227 0 PWM_CNTB[11]
rlabel metal2 23230 1588 23230 1588 0 PWM_CNTB[12]
rlabel metal2 29394 15249 29394 15249 0 PWM_CNTB[13]
rlabel metal2 29394 11033 29394 11033 0 PWM_CNTB[14]
rlabel metal1 9798 30294 9798 30294 0 PWM_CNTB[15]
rlabel metal1 11040 30226 11040 30226 0 PWM_CNTB[16]
rlabel metal2 29302 24667 29302 24667 0 PWM_CNTB[17]
rlabel metal3 751 4828 751 4828 0 PWM_CNTB[18]
rlabel metal2 7774 1588 7774 1588 0 PWM_CNTB[19]
rlabel metal2 29302 27149 29302 27149 0 PWM_CNTB[1]
rlabel metal3 29816 748 29816 748 0 PWM_CNTB[20]
rlabel metal1 16836 30226 16836 30226 0 PWM_CNTB[21]
rlabel metal3 751 23868 751 23868 0 PWM_CNTB[22]
rlabel metal1 7176 30226 7176 30226 0 PWM_CNTB[23]
rlabel metal1 12328 30226 12328 30226 0 PWM_CNTB[24]
rlabel metal2 29302 28883 29302 28883 0 PWM_CNTB[25]
rlabel metal3 29632 68 29632 68 0 PWM_CNTB[26]
rlabel metal1 14904 30226 14904 30226 0 PWM_CNTB[27]
rlabel metal2 11638 1554 11638 1554 0 PWM_CNTB[28]
rlabel metal2 29302 8347 29302 8347 0 PWM_CNTB[29]
rlabel metal2 29302 21029 29302 21029 0 PWM_CNTB[2]
rlabel metal3 751 16388 751 16388 0 PWM_CNTB[30]
rlabel metal1 18124 30226 18124 30226 0 PWM_CNTB[31]
rlabel metal2 5290 30719 5290 30719 0 PWM_CNTB[3]
rlabel metal2 24518 1588 24518 1588 0 PWM_CNTB[4]
rlabel metal3 751 3468 751 3468 0 PWM_CNTB[5]
rlabel metal2 20010 1588 20010 1588 0 PWM_CNTB[6]
rlabel metal2 1978 1588 1978 1588 0 PWM_CNTB[7]
rlabel metal2 9062 1588 9062 1588 0 PWM_CNTB[8]
rlabel metal2 29670 1588 29670 1588 0 PWM_CNTB[9]
rlabel metal3 751 748 751 748 0 PWM_OUTA
rlabel metal2 29394 9503 29394 9503 0 PWM_OUTB
rlabel metal2 22586 1588 22586 1588 0 TIMER_TOP[0]
rlabel metal3 1096 25908 1096 25908 0 TIMER_TOP[10]
rlabel via2 29302 3451 29302 3451 0 TIMER_TOP[11]
rlabel metal3 751 7548 751 7548 0 TIMER_TOP[12]
rlabel metal2 29302 13787 29302 13787 0 TIMER_TOP[13]
rlabel metal3 29770 22508 29770 22508 0 TIMER_TOP[14]
rlabel metal2 25806 1554 25806 1554 0 TIMER_TOP[15]
rlabel metal2 29302 23817 29302 23817 0 TIMER_TOP[16]
rlabel metal2 15502 1554 15502 1554 0 TIMER_TOP[17]
rlabel metal3 820 32708 820 32708 0 TIMER_TOP[18]
rlabel metal3 1050 13668 1050 13668 0 TIMER_TOP[19]
rlabel metal2 46 1554 46 1554 0 TIMER_TOP[1]
rlabel metal2 18722 1554 18722 1554 0 TIMER_TOP[20]
rlabel metal1 3956 30226 3956 30226 0 TIMER_TOP[21]
rlabel metal1 13708 30226 13708 30226 0 TIMER_TOP[22]
rlabel metal3 1050 8228 1050 8228 0 TIMER_TOP[23]
rlabel metal3 958 31348 958 31348 0 TIMER_TOP[24]
rlabel metal2 4554 1554 4554 1554 0 TIMER_TOP[25]
rlabel metal1 1426 2958 1426 2958 0 TIMER_TOP[26]
rlabel metal1 27922 30294 27922 30294 0 TIMER_TOP[27]
rlabel metal1 20792 30294 20792 30294 0 TIMER_TOP[28]
rlabel metal2 14214 1554 14214 1554 0 TIMER_TOP[29]
rlabel metal1 28474 30260 28474 30260 0 TIMER_TOP[2]
rlabel metal2 29302 5015 29302 5015 0 TIMER_TOP[30]
rlabel metal2 46 31256 46 31256 0 TIMER_TOP[31]
rlabel metal3 751 12308 751 12308 0 TIMER_TOP[3]
rlabel metal2 5842 1588 5842 1588 0 TIMER_TOP[4]
rlabel metal2 10350 1588 10350 1588 0 TIMER_TOP[5]
rlabel metal2 16146 1588 16146 1588 0 TIMER_TOP[6]
rlabel metal2 29302 19601 29302 19601 0 TIMER_TOP[7]
rlabel metal2 17434 1588 17434 1588 0 TIMER_TOP[8]
rlabel metal1 23920 30226 23920 30226 0 TIMER_TOP[9]
rlabel metal1 22632 30226 22632 30226 0 TMR_MODE[0]
rlabel metal1 1886 30294 1886 30294 0 TMR_MODE[1]
rlabel metal2 23782 4318 23782 4318 0 _0000_
rlabel metal1 14818 10234 14818 10234 0 _0001_
rlabel metal1 14848 11322 14848 11322 0 _0002_
rlabel metal1 14766 12410 14766 12410 0 _0003_
rlabel metal1 5290 12750 5290 12750 0 _0004_
rlabel metal1 7130 14314 7130 14314 0 _0005_
rlabel metal1 4554 13804 4554 13804 0 _0006_
rlabel metal1 3680 22202 3680 22202 0 _0007_
rlabel metal1 3075 24378 3075 24378 0 _0008_
rlabel metal1 4094 25466 4094 25466 0 _0009_
rlabel metal1 5888 27098 5888 27098 0 _0010_
rlabel metal2 23598 2788 23598 2788 0 _0011_
rlabel metal2 8142 27166 8142 27166 0 _0012_
rlabel metal2 8050 28254 8050 28254 0 _0013_
rlabel metal2 10534 28322 10534 28322 0 _0014_
rlabel metal1 11638 27336 11638 27336 0 _0015_
rlabel metal2 12926 28254 12926 28254 0 _0016_
rlabel metal2 14582 28560 14582 28560 0 _0017_
rlabel metal1 17296 27982 17296 27982 0 _0018_
rlabel metal2 18078 28356 18078 28356 0 _0019_
rlabel metal1 20148 28186 20148 28186 0 _0020_
rlabel metal1 20286 27370 20286 27370 0 _0021_
rlabel metal2 21298 3298 21298 3298 0 _0022_
rlabel metal2 23322 26214 23322 26214 0 _0023_
rlabel metal1 19872 25806 19872 25806 0 _0024_
rlabel metal1 19872 3638 19872 3638 0 _0025_
rlabel metal1 19872 3094 19872 3094 0 _0026_
rlabel metal1 18032 3094 18032 3094 0 _0027_
rlabel metal2 14674 3774 14674 3774 0 _0028_
rlabel metal2 13294 3400 13294 3400 0 _0029_
rlabel metal1 11270 3400 11270 3400 0 _0030_
rlabel metal1 10028 4046 10028 4046 0 _0031_
rlabel metal1 20874 22202 20874 22202 0 _0032_
rlabel metal2 20470 22746 20470 22746 0 _0033_
rlabel via1 23690 24106 23690 24106 0 _0034_
rlabel metal1 14444 14586 14444 14586 0 _0035_
rlabel metal1 21206 20026 21206 20026 0 _0036_
rlabel metal1 22034 20502 22034 20502 0 _0037_
rlabel metal2 25346 10846 25346 10846 0 _0038_
rlabel metal1 25576 16218 25576 16218 0 _0039_
rlabel metal2 25530 17816 25530 17816 0 _0040_
rlabel metal2 27738 17374 27738 17374 0 _0041_
rlabel metal2 27922 18462 27922 18462 0 _0042_
rlabel metal2 27922 20060 27922 20060 0 _0043_
rlabel metal2 25162 19618 25162 19618 0 _0044_
rlabel metal2 25346 21080 25346 21080 0 _0045_
rlabel metal1 25106 22202 25106 22202 0 _0046_
rlabel metal1 27646 21454 27646 21454 0 _0047_
rlabel metal2 27922 22814 27922 22814 0 _0048_
rlabel metal1 26818 9622 26818 9622 0 _0049_
rlabel metal2 28198 23970 28198 23970 0 _0050_
rlabel metal1 26036 23834 26036 23834 0 _0051_
rlabel metal2 28014 25636 28014 25636 0 _0052_
rlabel metal1 27830 27098 27830 27098 0 _0053_
rlabel metal1 25392 26010 25392 26010 0 _0054_
rlabel metal1 27462 27982 27462 27982 0 _0055_
rlabel metal1 25208 27642 25208 27642 0 _0056_
rlabel metal1 23322 28594 23322 28594 0 _0057_
rlabel metal1 23745 27642 23745 27642 0 _0058_
rlabel metal1 24518 26554 24518 26554 0 _0059_
rlabel metal1 27968 10098 27968 10098 0 _0060_
rlabel metal2 24242 24548 24242 24548 0 _0061_
rlabel metal1 22908 24378 22908 24378 0 _0062_
rlabel metal1 27692 11798 27692 11798 0 _0063_
rlabel metal2 25714 12444 25714 12444 0 _0064_
rlabel metal1 25024 12954 25024 12954 0 _0065_
rlabel metal2 27922 13532 27922 13532 0 _0066_
rlabel metal1 28099 14586 28099 14586 0 _0067_
rlabel metal1 27646 15946 27646 15946 0 _0068_
rlabel metal1 25300 14314 25300 14314 0 _0069_
rlabel metal2 23506 13736 23506 13736 0 _0070_
rlabel metal1 25445 11798 25445 11798 0 _0071_
rlabel metal2 21942 13090 21942 13090 0 _0072_
rlabel metal2 24150 10472 24150 10472 0 _0073_
rlabel metal1 20339 12886 20339 12886 0 _0074_
rlabel metal2 17710 13022 17710 13022 0 _0075_
rlabel metal2 20102 8738 20102 8738 0 _0076_
rlabel metal1 15548 8058 15548 8058 0 _0077_
rlabel metal1 8747 8874 8747 8874 0 _0078_
rlabel metal1 8103 5270 8103 5270 0 _0079_
rlabel metal2 2438 6562 2438 6562 0 _0080_
rlabel metal1 5612 5338 5612 5338 0 _0081_
rlabel metal1 5198 8602 5198 8602 0 _0082_
rlabel metal2 2162 9384 2162 9384 0 _0083_
rlabel metal2 2162 13022 2162 13022 0 _0084_
rlabel metal2 3450 14110 3450 14110 0 _0085_
rlabel metal2 2622 15912 2622 15912 0 _0086_
rlabel metal2 2806 19142 2806 19142 0 _0087_
rlabel metal1 4002 21114 4002 21114 0 _0088_
rlabel metal1 4692 20026 4692 20026 0 _0089_
rlabel metal1 6893 16150 6893 16150 0 _0090_
rlabel metal1 13577 18326 13577 18326 0 _0091_
rlabel metal2 14306 16286 14306 16286 0 _0092_
rlabel metal2 6946 17442 6946 17442 0 _0093_
rlabel metal1 16468 16966 16468 16966 0 _0094_
rlabel metal1 20056 17306 20056 17306 0 _0095_
rlabel metal1 16659 13226 16659 13226 0 _0096_
rlabel metal1 20976 14042 20976 14042 0 _0097_
rlabel metal1 24472 15334 24472 15334 0 _0098_
rlabel metal1 24663 19414 24663 19414 0 _0099_
rlabel metal1 24564 17850 24564 17850 0 _0100_
rlabel metal2 24058 16286 24058 16286 0 _0101_
rlabel metal2 25070 22780 25070 22780 0 _0102_
rlabel metal1 26266 11016 26266 11016 0 _0103_
rlabel metal2 27370 9384 27370 9384 0 _0104_
rlabel metal2 29026 9826 29026 9826 0 _0105_
rlabel metal1 28934 11322 28934 11322 0 _0106_
rlabel metal1 27147 12138 27147 12138 0 _0107_
rlabel metal1 26220 13498 26220 13498 0 _0108_
rlabel metal1 28888 12954 28888 12954 0 _0109_
rlabel metal2 28934 14178 28934 14178 0 _0110_
rlabel metal2 28934 16286 28934 16286 0 _0111_
rlabel metal2 26266 14586 26266 14586 0 _0112_
rlabel metal1 26358 16218 26358 16218 0 _0113_
rlabel metal1 26312 18054 26312 18054 0 _0114_
rlabel metal1 28704 16762 28704 16762 0 _0115_
rlabel metal1 28888 17850 28888 17850 0 _0116_
rlabel metal2 28934 19618 28934 19618 0 _0117_
rlabel metal2 25990 19618 25990 19618 0 _0118_
rlabel metal1 26266 20570 26266 20570 0 _0119_
rlabel metal1 26641 21930 26641 21930 0 _0120_
rlabel metal1 28796 21114 28796 21114 0 _0121_
rlabel metal2 28934 22372 28934 22372 0 _0122_
rlabel metal2 28934 23970 28934 23970 0 _0123_
rlabel metal2 26358 24344 26358 24344 0 _0124_
rlabel metal1 28934 25466 28934 25466 0 _0125_
rlabel metal2 28934 27234 28934 27234 0 _0126_
rlabel metal1 26220 26010 26220 26010 0 _0127_
rlabel metal1 28803 28458 28803 28458 0 _0128_
rlabel metal1 26503 28118 26503 28118 0 _0129_
rlabel metal1 23368 29002 23368 29002 0 _0130_
rlabel metal1 22632 27098 22632 27098 0 _0131_
rlabel metal1 24656 26010 24656 26010 0 _0132_
rlabel metal1 25208 24378 25208 24378 0 _0133_
rlabel metal1 22540 24378 22540 24378 0 _0134_
rlabel metal1 22073 22678 22073 22678 0 _0135_
rlabel metal1 22639 21930 22639 21930 0 _0136_
rlabel metal2 24518 4318 24518 4318 0 _0137_
rlabel metal1 25031 3094 25031 3094 0 _0138_
rlabel metal1 21988 3162 21988 3162 0 _0139_
rlabel metal2 20470 4318 20470 4318 0 _0140_
rlabel metal2 19366 2720 19366 2720 0 _0141_
rlabel metal2 17066 2822 17066 2822 0 _0142_
rlabel metal1 15456 3162 15456 3162 0 _0143_
rlabel metal1 14727 3094 14727 3094 0 _0144_
rlabel metal1 12052 3162 12052 3162 0 _0145_
rlabel metal2 9982 3944 9982 3944 0 _0146_
rlabel metal2 14950 9792 14950 9792 0 _0147_
rlabel metal1 16383 11050 16383 11050 0 _0148_
rlabel metal1 15824 12410 15824 12410 0 _0149_
rlabel metal1 5428 12410 5428 12410 0 _0150_
rlabel metal1 8793 14314 8793 14314 0 _0151_
rlabel metal2 5474 14178 5474 14178 0 _0152_
rlabel metal1 4002 22066 4002 22066 0 _0153_
rlabel metal2 3266 24004 3266 24004 0 _0154_
rlabel metal2 4738 26078 4738 26078 0 _0155_
rlabel metal1 5888 27846 5888 27846 0 _0156_
rlabel metal1 9108 27302 9108 27302 0 _0157_
rlabel metal2 9062 28254 9062 28254 0 _0158_
rlabel metal1 11224 29002 11224 29002 0 _0159_
rlabel metal1 12558 27098 12558 27098 0 _0160_
rlabel metal2 13662 28254 13662 28254 0 _0161_
rlabel metal1 15732 28730 15732 28730 0 _0162_
rlabel metal1 17112 27574 17112 27574 0 _0163_
rlabel metal1 18860 28730 18860 28730 0 _0164_
rlabel metal1 21252 28186 21252 28186 0 _0165_
rlabel metal1 21252 27098 21252 27098 0 _0166_
rlabel metal2 22310 25704 22310 25704 0 _0167_
rlabel metal2 21482 25704 21482 25704 0 _0168_
rlabel metal1 24479 20502 24479 20502 0 _0169_
rlabel metal1 22540 20570 22540 20570 0 _0170_
rlabel metal2 16238 14824 16238 14824 0 _0171_
rlabel metal1 22622 13702 22622 13702 0 _0172_
rlabel metal2 23966 11866 23966 11866 0 _0173_
rlabel metal2 20930 13090 20930 13090 0 _0174_
rlabel metal1 23000 10234 23000 10234 0 _0175_
rlabel metal1 19090 12410 19090 12410 0 _0176_
rlabel metal1 17112 12410 17112 12410 0 _0177_
rlabel metal1 19688 8602 19688 8602 0 _0178_
rlabel metal2 14766 8670 14766 8670 0 _0179_
rlabel metal1 7084 8602 7084 8602 0 _0180_
rlabel metal2 6670 5406 6670 5406 0 _0181_
rlabel via1 1695 6970 1695 6970 0 _0182_
rlabel metal1 4600 5338 4600 5338 0 _0183_
rlabel metal1 4462 9010 4462 9010 0 _0184_
rlabel metal2 2346 9316 2346 9316 0 _0185_
rlabel metal1 1794 12410 1794 12410 0 _0186_
rlabel metal2 3818 13600 3818 13600 0 _0187_
rlabel metal1 3266 15980 3266 15980 0 _0188_
rlabel metal2 1702 19550 1702 19550 0 _0189_
rlabel metal1 3496 18938 3496 18938 0 _0190_
rlabel metal1 4738 19278 4738 19278 0 _0191_
rlabel metal1 6624 15674 6624 15674 0 _0192_
rlabel metal1 11960 17850 11960 17850 0 _0193_
rlabel metal2 13570 16286 13570 16286 0 _0194_
rlabel metal2 7130 17408 7130 17408 0 _0195_
rlabel metal1 15548 16218 15548 16218 0 _0196_
rlabel metal2 19734 17408 19734 17408 0 _0197_
rlabel metal1 15502 13362 15502 13362 0 _0198_
rlabel metal1 19918 14042 19918 14042 0 _0199_
rlabel metal1 23276 15062 23276 15062 0 _0200_
rlabel metal2 22494 19108 22494 19108 0 _0201_
rlabel metal1 23230 18156 23230 18156 0 _0202_
rlabel metal2 24518 16422 24518 16422 0 _0203_
rlabel metal2 11638 12274 11638 12274 0 _0204_
rlabel metal1 11960 13498 11960 13498 0 _0205_
rlabel metal1 12512 13430 12512 13430 0 _0206_
rlabel metal1 12156 13974 12156 13974 0 _0207_
rlabel metal2 12190 15963 12190 15963 0 _0208_
rlabel metal2 12466 23596 12466 23596 0 _0209_
rlabel metal2 11086 23290 11086 23290 0 _0210_
rlabel metal1 11822 23018 11822 23018 0 _0211_
rlabel metal1 13340 23222 13340 23222 0 _0212_
rlabel metal1 16560 22746 16560 22746 0 _0213_
rlabel metal1 16652 23290 16652 23290 0 _0214_
rlabel metal1 18170 23120 18170 23120 0 _0215_
rlabel metal1 15180 23086 15180 23086 0 _0216_
rlabel metal1 15870 23290 15870 23290 0 _0217_
rlabel metal2 18078 22916 18078 22916 0 _0218_
rlabel metal1 16836 22474 16836 22474 0 _0219_
rlabel metal2 16882 22848 16882 22848 0 _0220_
rlabel metal1 15272 23018 15272 23018 0 _0221_
rlabel metal2 15134 23290 15134 23290 0 _0222_
rlabel metal2 17986 23460 17986 23460 0 _0223_
rlabel metal1 16790 23052 16790 23052 0 _0224_
rlabel metal1 17342 23120 17342 23120 0 _0225_
rlabel metal1 18814 23154 18814 23154 0 _0226_
rlabel metal1 17802 23052 17802 23052 0 _0227_
rlabel metal2 10166 12002 10166 12002 0 _0228_
rlabel metal1 10166 12886 10166 12886 0 _0229_
rlabel metal1 9476 12954 9476 12954 0 _0230_
rlabel metal1 10166 13702 10166 13702 0 _0231_
rlabel metal2 10534 12036 10534 12036 0 _0232_
rlabel metal2 10074 12512 10074 12512 0 _0233_
rlabel metal2 22586 6086 22586 6086 0 _0234_
rlabel metal1 23322 6221 23322 6221 0 _0235_
rlabel metal1 22126 6256 22126 6256 0 _0236_
rlabel metal1 20700 6290 20700 6290 0 _0237_
rlabel metal2 18262 5882 18262 5882 0 _0238_
rlabel metal1 18078 5610 18078 5610 0 _0239_
rlabel metal1 18400 5678 18400 5678 0 _0240_
rlabel metal1 14582 5712 14582 5712 0 _0241_
rlabel metal1 14812 5338 14812 5338 0 _0242_
rlabel metal1 13294 5338 13294 5338 0 _0243_
rlabel metal1 11914 5712 11914 5712 0 _0244_
rlabel metal1 11776 5338 11776 5338 0 _0245_
rlabel metal2 11730 5882 11730 5882 0 _0246_
rlabel metal2 11546 6630 11546 6630 0 _0247_
rlabel metal1 11914 7514 11914 7514 0 _0248_
rlabel metal1 11132 11866 11132 11866 0 _0249_
rlabel metal1 9890 12240 9890 12240 0 _0250_
rlabel metal2 8832 17204 8832 17204 0 _0251_
rlabel metal1 7728 24786 7728 24786 0 _0252_
rlabel metal1 6118 26010 6118 26010 0 _0253_
rlabel metal2 7590 25568 7590 25568 0 _0254_
rlabel metal2 5382 24582 5382 24582 0 _0255_
rlabel metal2 5658 24106 5658 24106 0 _0256_
rlabel metal2 7038 25228 7038 25228 0 _0257_
rlabel metal1 7038 24786 7038 24786 0 _0258_
rlabel metal2 5934 24548 5934 24548 0 _0259_
rlabel metal1 9246 24106 9246 24106 0 _0260_
rlabel metal1 9154 24140 9154 24140 0 _0261_
rlabel metal1 5382 24650 5382 24650 0 _0262_
rlabel metal1 6394 25874 6394 25874 0 _0263_
rlabel metal2 7682 25466 7682 25466 0 _0264_
rlabel metal1 7590 24854 7590 24854 0 _0265_
rlabel metal2 8970 24378 8970 24378 0 _0266_
rlabel metal2 14490 24004 14490 24004 0 _0267_
rlabel metal2 20010 23154 20010 23154 0 _0268_
rlabel metal1 21068 23494 21068 23494 0 _0269_
rlabel via1 20930 23698 20930 23698 0 _0270_
rlabel metal1 17756 23494 17756 23494 0 _0271_
rlabel metal1 18814 23596 18814 23596 0 _0272_
rlabel metal1 21068 24242 21068 24242 0 _0273_
rlabel metal1 19044 24038 19044 24038 0 _0274_
rlabel metal1 18584 24174 18584 24174 0 _0275_
rlabel metal2 18446 24242 18446 24242 0 _0276_
rlabel metal1 18308 23766 18308 23766 0 _0277_
rlabel metal2 19826 23052 19826 23052 0 _0278_
rlabel metal2 19642 24140 19642 24140 0 _0279_
rlabel metal2 19918 23902 19918 23902 0 _0280_
rlabel metal1 20010 22542 20010 22542 0 _0281_
rlabel metal1 10626 10438 10626 10438 0 _0282_
rlabel metal2 10626 11526 10626 11526 0 _0283_
rlabel metal2 17250 6494 17250 6494 0 _0284_
rlabel metal1 24288 7718 24288 7718 0 _0285_
rlabel metal1 24426 7514 24426 7514 0 _0286_
rlabel metal1 23966 7786 23966 7786 0 _0287_
rlabel metal1 19734 7888 19734 7888 0 _0288_
rlabel metal2 20102 7684 20102 7684 0 _0289_
rlabel metal1 19320 6630 19320 6630 0 _0290_
rlabel metal1 18446 6290 18446 6290 0 _0291_
rlabel metal2 17066 5542 17066 5542 0 _0292_
rlabel metal1 11500 5202 11500 5202 0 _0293_
rlabel metal2 11086 5508 11086 5508 0 _0294_
rlabel metal1 10672 5270 10672 5270 0 _0295_
rlabel metal1 10626 5202 10626 5202 0 _0296_
rlabel metal2 10258 5644 10258 5644 0 _0297_
rlabel metal1 10028 5338 10028 5338 0 _0298_
rlabel metal2 10994 8126 10994 8126 0 _0299_
rlabel metal2 10166 9690 10166 9690 0 _0300_
rlabel metal1 10120 9690 10120 9690 0 _0301_
rlabel metal1 10120 10234 10120 10234 0 _0302_
rlabel metal2 11132 13702 11132 13702 0 _0303_
rlabel metal1 11960 20774 11960 20774 0 _0304_
rlabel metal2 9430 20944 9430 20944 0 _0305_
rlabel metal1 9384 20570 9384 20570 0 _0306_
rlabel metal2 9982 21284 9982 21284 0 _0307_
rlabel metal1 12742 21930 12742 21930 0 _0308_
rlabel metal2 11270 21930 11270 21930 0 _0309_
rlabel metal2 8418 21726 8418 21726 0 _0310_
rlabel metal2 7406 21658 7406 21658 0 _0311_
rlabel via1 12573 21998 12573 21998 0 _0312_
rlabel metal1 8234 21488 8234 21488 0 _0313_
rlabel metal1 8602 21624 8602 21624 0 _0314_
rlabel metal2 11914 21114 11914 21114 0 _0315_
rlabel metal1 11960 22066 11960 22066 0 _0316_
rlabel metal1 8188 21930 8188 21930 0 _0317_
rlabel metal1 8786 21998 8786 21998 0 _0318_
rlabel metal2 9614 21692 9614 21692 0 _0319_
rlabel metal1 9890 21658 9890 21658 0 _0320_
rlabel metal1 12098 20910 12098 20910 0 _0321_
rlabel metal1 16330 20400 16330 20400 0 _0322_
rlabel metal1 17710 19788 17710 19788 0 _0323_
rlabel metal2 15594 21284 15594 21284 0 _0324_
rlabel metal2 18078 20196 18078 20196 0 _0325_
rlabel metal2 18170 19380 18170 19380 0 _0326_
rlabel metal1 16652 20230 16652 20230 0 _0327_
rlabel metal2 16606 21114 16606 21114 0 _0328_
rlabel metal1 16974 21590 16974 21590 0 _0329_
rlabel metal2 17066 21148 17066 21148 0 _0330_
rlabel metal2 16882 20604 16882 20604 0 _0331_
rlabel metal1 14490 20502 14490 20502 0 _0332_
rlabel metal1 16054 20536 16054 20536 0 _0333_
rlabel metal1 17618 20434 17618 20434 0 _0334_
rlabel metal1 16698 20366 16698 20366 0 _0335_
rlabel metal2 16698 20604 16698 20604 0 _0336_
rlabel metal2 17894 20026 17894 20026 0 _0337_
rlabel metal1 18262 20026 18262 20026 0 _0338_
rlabel metal1 20148 19482 20148 19482 0 _0339_
rlabel metal1 17894 19686 17894 19686 0 _0340_
rlabel metal1 21298 19482 21298 19482 0 _0341_
rlabel metal2 21206 20706 21206 20706 0 _0342_
rlabel via1 19550 20434 19550 20434 0 _0343_
rlabel metal1 19274 20468 19274 20468 0 _0344_
rlabel metal1 19274 20570 19274 20570 0 _0345_
rlabel metal1 21022 20944 21022 20944 0 _0346_
rlabel metal2 21022 20060 21022 20060 0 _0347_
rlabel metal1 20795 19482 20795 19482 0 _0348_
rlabel metal2 8694 19006 8694 19006 0 _0349_
rlabel metal2 8786 19584 8786 19584 0 _0350_
rlabel metal1 6946 19380 6946 19380 0 _0351_
rlabel metal2 5658 19618 5658 19618 0 _0352_
rlabel metal2 6854 20740 6854 20740 0 _0353_
rlabel metal2 6578 20298 6578 20298 0 _0354_
rlabel metal2 6578 21148 6578 21148 0 _0355_
rlabel metal1 6026 20264 6026 20264 0 _0356_
rlabel metal2 6394 20026 6394 20026 0 _0357_
rlabel metal2 7038 19516 7038 19516 0 _0358_
rlabel metal1 7222 18666 7222 18666 0 _0359_
rlabel metal1 6486 21964 6486 21964 0 _0360_
rlabel metal2 7498 19686 7498 19686 0 _0361_
rlabel metal2 20562 8058 20562 8058 0 _0362_
rlabel metal2 23414 9146 23414 9146 0 _0363_
rlabel metal1 23460 8602 23460 8602 0 _0364_
rlabel metal1 23690 8908 23690 8908 0 _0365_
rlabel metal1 21390 7888 21390 7888 0 _0366_
rlabel metal1 18584 6698 18584 6698 0 _0367_
rlabel metal1 17940 6766 17940 6766 0 _0368_
rlabel metal2 17526 6970 17526 6970 0 _0369_
rlabel metal1 15870 6358 15870 6358 0 _0370_
rlabel metal2 8786 5950 8786 5950 0 _0371_
rlabel metal1 8832 5814 8832 5814 0 _0372_
rlabel metal1 8648 5338 8648 5338 0 _0373_
rlabel metal2 8326 6324 8326 6324 0 _0374_
rlabel metal1 8188 6426 8188 6426 0 _0375_
rlabel metal1 8694 7310 8694 7310 0 _0376_
rlabel metal1 8004 6970 8004 6970 0 _0377_
rlabel metal1 8786 6970 8786 6970 0 _0378_
rlabel metal1 8050 6800 8050 6800 0 _0379_
rlabel metal2 7866 8432 7866 8432 0 _0380_
rlabel metal2 8326 11968 8326 11968 0 _0381_
rlabel metal2 7590 12988 7590 12988 0 _0382_
rlabel metal1 7544 12614 7544 12614 0 _0383_
rlabel metal1 7958 12614 7958 12614 0 _0384_
rlabel metal1 9200 10642 9200 10642 0 _0385_
rlabel metal1 9154 10438 9154 10438 0 _0386_
rlabel metal1 8418 10030 8418 10030 0 _0387_
rlabel metal2 7682 10948 7682 10948 0 _0388_
rlabel metal1 7958 10778 7958 10778 0 _0389_
rlabel via1 7878 11798 7878 11798 0 _0390_
rlabel metal1 7958 19822 7958 19822 0 _0391_
rlabel metal2 7222 19652 7222 19652 0 _0392_
rlabel metal2 7130 21182 7130 21182 0 _0393_
rlabel metal1 7682 19856 7682 19856 0 _0394_
rlabel via2 7958 19669 7958 19669 0 _0395_
rlabel metal1 15318 19924 15318 19924 0 _0396_
rlabel metal2 20240 20434 20240 20434 0 _0397_
rlabel metal2 20654 19958 20654 19958 0 _0398_
rlabel metal2 19826 20094 19826 20094 0 _0399_
rlabel metal1 20378 19788 20378 19788 0 _0400_
rlabel metal1 27968 10642 27968 10642 0 _0401_
rlabel metal1 27830 11322 27830 11322 0 _0402_
rlabel metal1 25898 12852 25898 12852 0 _0403_
rlabel metal2 27554 13362 27554 13362 0 _0404_
rlabel metal1 27646 14586 27646 14586 0 _0405_
rlabel metal1 26312 14858 26312 14858 0 _0406_
rlabel metal2 25438 16524 25438 16524 0 _0407_
rlabel metal1 27508 16762 27508 16762 0 _0408_
rlabel metal1 28014 18768 28014 18768 0 _0409_
rlabel metal1 26082 19210 26082 19210 0 _0410_
rlabel metal1 26036 21522 26036 21522 0 _0411_
rlabel metal1 27416 21114 27416 21114 0 _0412_
rlabel metal1 27968 23086 27968 23086 0 _0413_
rlabel metal1 26772 23562 26772 23562 0 _0414_
rlabel metal1 27784 25262 27784 25262 0 _0415_
rlabel metal1 26266 25738 26266 25738 0 _0416_
rlabel metal2 25346 28050 25346 28050 0 _0417_
rlabel metal2 24518 28356 24518 28356 0 _0418_
rlabel metal1 23782 26350 23782 26350 0 _0419_
rlabel metal2 23138 24718 23138 24718 0 _0420_
rlabel metal1 17572 17646 17572 17646 0 _0421_
rlabel metal1 21206 18938 21206 18938 0 _0422_
rlabel metal1 18538 18836 18538 18836 0 _0423_
rlabel metal1 17204 20434 17204 20434 0 _0424_
rlabel metal2 17342 18785 17342 18785 0 _0425_
rlabel metal1 19734 21386 19734 21386 0 _0426_
rlabel metal2 15042 19550 15042 19550 0 _0427_
rlabel metal2 14582 19006 14582 19006 0 _0428_
rlabel metal2 8418 19040 8418 19040 0 _0429_
rlabel metal1 7268 22066 7268 22066 0 _0430_
rlabel metal1 11039 21998 11039 21998 0 _0431_
rlabel metal1 9614 18734 9614 18734 0 _0432_
rlabel metal1 9016 20026 9016 20026 0 _0433_
rlabel metal2 6210 20434 6210 20434 0 _0434_
rlabel via1 6485 20910 6485 20910 0 _0435_
rlabel metal2 8418 20604 8418 20604 0 _0436_
rlabel metal2 13570 20604 13570 20604 0 _0437_
rlabel metal1 7774 12784 7774 12784 0 _0438_
rlabel metal1 8970 9690 8970 9690 0 _0439_
rlabel metal1 8970 7412 8970 7412 0 _0440_
rlabel metal1 8786 7378 8786 7378 0 _0441_
rlabel metal1 8648 6290 8648 6290 0 _0442_
rlabel metal2 9614 6528 9614 6528 0 _0443_
rlabel metal1 12604 8466 12604 8466 0 _0444_
rlabel metal1 15594 6188 15594 6188 0 _0445_
rlabel metal1 17480 10710 17480 10710 0 _0446_
rlabel metal2 20102 10404 20102 10404 0 _0447_
rlabel metal1 21068 8806 21068 8806 0 _0448_
rlabel metal1 23966 8432 23966 8432 0 _0449_
rlabel via1 23690 8483 23690 8483 0 _0450_
rlabel metal2 24150 9078 24150 9078 0 _0451_
rlabel metal2 18722 26656 18722 26656 0 _0452_
rlabel metal1 18446 25908 18446 25908 0 _0453_
rlabel metal2 18170 26078 18170 26078 0 _0454_
rlabel metal1 17342 26384 17342 26384 0 _0455_
rlabel metal1 16836 20026 16836 20026 0 _0456_
rlabel metal1 16882 19380 16882 19380 0 _0457_
rlabel metal1 14674 24582 14674 24582 0 _0458_
rlabel metal1 12972 21114 12972 21114 0 _0459_
rlabel metal2 13432 22066 13432 22066 0 _0460_
rlabel metal1 12788 22066 12788 22066 0 _0461_
rlabel metal2 11730 20060 11730 20060 0 _0462_
rlabel metal1 14076 13974 14076 13974 0 _0463_
rlabel metal1 12190 9554 12190 9554 0 _0464_
rlabel metal1 12098 9962 12098 9962 0 _0465_
rlabel metal2 13110 7174 13110 7174 0 _0466_
rlabel via1 16790 6834 16790 6834 0 _0467_
rlabel via1 21022 5542 21022 5542 0 _0468_
rlabel metal2 21298 7956 21298 7956 0 _0469_
rlabel metal1 19964 13498 19964 13498 0 _0470_
rlabel metal1 20102 21930 20102 21930 0 _0471_
rlabel metal1 19642 22610 19642 22610 0 _0472_
rlabel metal1 19826 24650 19826 24650 0 _0473_
rlabel metal1 17711 22576 17711 22576 0 _0474_
rlabel metal2 17434 24599 17434 24599 0 _0475_
rlabel metal1 18446 24106 18446 24106 0 _0476_
rlabel metal1 15042 23766 15042 23766 0 _0477_
rlabel metal2 14490 25568 14490 25568 0 _0478_
rlabel metal2 8694 24446 8694 24446 0 _0479_
rlabel via1 9982 24378 9982 24378 0 _0480_
rlabel metal1 9200 25126 9200 25126 0 _0481_
rlabel metal2 10350 26622 10350 26622 0 _0482_
rlabel metal1 6348 25806 6348 25806 0 _0483_
rlabel metal1 10212 25262 10212 25262 0 _0484_
rlabel metal1 10902 25262 10902 25262 0 _0485_
rlabel via1 7756 25874 7756 25874 0 _0486_
rlabel metal1 7498 13702 7498 13702 0 _0487_
rlabel metal2 9246 14178 9246 14178 0 _0488_
rlabel metal1 13386 11696 13386 11696 0 _0489_
rlabel metal1 14444 7446 14444 7446 0 _0490_
rlabel metal2 11822 7616 11822 7616 0 _0491_
rlabel metal2 13754 6800 13754 6800 0 _0492_
rlabel viali 11822 5205 11822 5205 0 _0493_
rlabel metal2 15502 5508 15502 5508 0 _0494_
rlabel metal2 17480 5202 17480 5202 0 _0495_
rlabel metal2 19090 5372 19090 5372 0 _0496_
rlabel metal2 19274 5542 19274 5542 0 _0497_
rlabel viali 20511 6290 20511 6290 0 _0498_
rlabel metal1 23368 3706 23368 3706 0 _0499_
rlabel metal1 23598 6154 23598 6154 0 _0500_
rlabel metal1 24150 6358 24150 6358 0 _0501_
rlabel metal1 17158 22202 17158 22202 0 _0502_
rlabel metal1 15134 21522 15134 21522 0 _0503_
rlabel metal1 14582 21590 14582 21590 0 _0504_
rlabel metal1 12834 22542 12834 22542 0 _0505_
rlabel metal1 12972 23290 12972 23290 0 _0506_
rlabel metal1 9798 22746 9798 22746 0 _0507_
rlabel metal2 9338 21590 9338 21590 0 _0508_
rlabel metal1 8326 21386 8326 21386 0 _0509_
rlabel metal1 7728 23222 7728 23222 0 _0510_
rlabel metal1 7981 23086 7981 23086 0 _0511_
rlabel metal2 7774 22542 7774 22542 0 _0512_
rlabel metal2 10166 14586 10166 14586 0 _0513_
rlabel metal2 10902 13770 10902 13770 0 _0514_
rlabel metal1 10856 11254 10856 11254 0 _0515_
rlabel metal1 10534 9996 10534 9996 0 _0516_
rlabel metal1 11776 9486 11776 9486 0 _0517_
rlabel metal2 13846 8262 13846 8262 0 _0518_
rlabel metal2 21114 6154 21114 6154 0 _0519_
rlabel metal2 22310 20519 22310 20519 0 _0520_
rlabel metal1 21344 20434 21344 20434 0 _0521_
rlabel metal1 21160 21658 21160 21658 0 _0522_
rlabel metal1 19366 21522 19366 21522 0 _0523_
rlabel metal2 15318 21760 15318 21760 0 _0524_
rlabel metal1 14720 22066 14720 22066 0 _0525_
rlabel metal1 8257 25874 8257 25874 0 _0526_
rlabel metal1 6902 21998 6902 21998 0 _0527_
rlabel metal1 6532 21522 6532 21522 0 _0528_
rlabel metal1 6394 21590 6394 21590 0 _0529_
rlabel metal1 5750 22576 5750 22576 0 _0530_
rlabel metal1 5842 22678 5842 22678 0 _0531_
rlabel metal1 8142 13192 8142 13192 0 _0532_
rlabel metal1 8142 12954 8142 12954 0 _0533_
rlabel metal1 8970 12818 8970 12818 0 _0534_
rlabel metal1 9430 11322 9430 11322 0 _0535_
rlabel metal2 7958 7548 7958 7548 0 _0536_
rlabel metal1 11086 19210 11086 19210 0 _0537_
rlabel metal2 13386 20876 13386 20876 0 _0538_
rlabel metal2 13064 20434 13064 20434 0 _0539_
rlabel metal1 11638 19924 11638 19924 0 _0540_
rlabel metal1 11914 19958 11914 19958 0 _0541_
rlabel metal1 10994 19856 10994 19856 0 _0542_
rlabel metal1 10442 19346 10442 19346 0 _0543_
rlabel metal1 10856 19754 10856 19754 0 _0544_
rlabel metal1 11178 19788 11178 19788 0 _0545_
rlabel metal2 10810 21114 10810 21114 0 _0546_
rlabel metal2 10994 19108 10994 19108 0 _0547_
rlabel metal1 10810 19482 10810 19482 0 _0548_
rlabel metal1 12581 19822 12581 19822 0 _0549_
rlabel metal1 13018 19346 13018 19346 0 _0550_
rlabel metal1 13202 15130 13202 15130 0 _0551_
rlabel metal1 9752 9010 9752 9010 0 _0552_
rlabel metal1 10810 8874 10810 8874 0 _0553_
rlabel metal1 22356 7514 22356 7514 0 _0554_
rlabel via1 22677 7854 22677 7854 0 _0555_
rlabel metal2 22770 7922 22770 7922 0 _0556_
rlabel metal1 21298 7480 21298 7480 0 _0557_
rlabel metal1 18814 6970 18814 6970 0 _0558_
rlabel metal2 21482 7582 21482 7582 0 _0559_
rlabel metal1 18630 7276 18630 7276 0 _0560_
rlabel metal1 19136 7310 19136 7310 0 _0561_
rlabel metal1 15686 7412 15686 7412 0 _0562_
rlabel metal1 15778 7276 15778 7276 0 _0563_
rlabel metal2 15318 7140 15318 7140 0 _0564_
rlabel metal1 15824 7514 15824 7514 0 _0565_
rlabel metal1 10212 7378 10212 7378 0 _0566_
rlabel metal2 10534 8092 10534 8092 0 _0567_
rlabel metal2 10350 8500 10350 8500 0 _0568_
rlabel metal1 11086 8908 11086 8908 0 _0569_
rlabel metal1 12745 8602 12745 8602 0 _0570_
rlabel metal1 12650 8976 12650 8976 0 _0571_
rlabel metal1 13478 9010 13478 9010 0 _0572_
rlabel viali 11178 8942 11178 8942 0 _0573_
rlabel metal1 12374 8908 12374 8908 0 _0574_
rlabel metal1 13846 8908 13846 8908 0 _0575_
rlabel metal1 13110 9044 13110 9044 0 _0576_
rlabel metal1 13156 15470 13156 15470 0 _0577_
rlabel metal1 12696 15130 12696 15130 0 _0578_
rlabel metal2 13294 17544 13294 17544 0 _0579_
rlabel metal1 13248 20570 13248 20570 0 _0580_
rlabel metal1 12591 20366 12591 20366 0 _0581_
rlabel metal1 12156 19346 12156 19346 0 _0582_
rlabel metal1 12328 19482 12328 19482 0 _0583_
rlabel via1 15213 18326 15213 18326 0 _0584_
rlabel metal2 17066 18428 17066 18428 0 _0585_
rlabel metal2 14398 19125 14398 19125 0 _0586_
rlabel metal1 15916 18190 15916 18190 0 _0587_
rlabel metal1 16698 18224 16698 18224 0 _0588_
rlabel metal2 15870 18938 15870 18938 0 _0589_
rlabel metal1 15686 18156 15686 18156 0 _0590_
rlabel metal1 14628 18802 14628 18802 0 _0591_
rlabel metal2 15318 18904 15318 18904 0 _0592_
rlabel metal2 17526 18564 17526 18564 0 _0593_
rlabel metal1 16146 18326 16146 18326 0 _0594_
rlabel metal2 15686 17850 15686 17850 0 _0595_
rlabel metal1 15502 18734 15502 18734 0 _0596_
rlabel via1 16790 18258 16790 18258 0 _0597_
rlabel metal1 16882 17714 16882 17714 0 _0598_
rlabel metal1 16146 17578 16146 17578 0 _0599_
rlabel metal1 15042 15504 15042 15504 0 _0600_
rlabel metal1 22724 11322 22724 11322 0 _0601_
rlabel metal2 21666 16762 21666 16762 0 _0602_
rlabel metal1 21160 15674 21160 15674 0 _0603_
rlabel metal2 18354 10132 18354 10132 0 _0604_
rlabel metal1 20470 16218 20470 16218 0 _0605_
rlabel metal1 13754 15436 13754 15436 0 _0606_
rlabel metal1 8970 17714 8970 17714 0 _0607_
rlabel metal1 9200 16218 9200 16218 0 _0608_
rlabel metal1 11086 17544 11086 17544 0 _0609_
rlabel metal1 12144 16218 12144 16218 0 _0610_
rlabel metal2 6578 8772 6578 8772 0 _0611_
rlabel metal2 5750 10404 5750 10404 0 _0612_
rlabel metal1 6716 10710 6716 10710 0 _0613_
rlabel metal1 7176 10778 7176 10778 0 _0614_
rlabel metal1 14352 15470 14352 15470 0 _0615_
rlabel metal1 17710 8398 17710 8398 0 _0616_
rlabel metal1 18998 11118 18998 11118 0 _0617_
rlabel metal1 19228 10778 19228 10778 0 _0618_
rlabel metal2 20010 11322 20010 11322 0 _0619_
rlabel metal1 21298 9520 21298 9520 0 _0620_
rlabel metal1 20148 10778 20148 10778 0 _0621_
rlabel metal1 21482 9588 21482 9588 0 _0622_
rlabel metal2 21298 10914 21298 10914 0 _0623_
rlabel metal2 22494 11696 22494 11696 0 _0624_
rlabel metal2 22310 11696 22310 11696 0 _0625_
rlabel metal1 22770 12274 22770 12274 0 _0626_
rlabel metal1 21436 10982 21436 10982 0 _0627_
rlabel metal1 21758 10778 21758 10778 0 _0628_
rlabel metal2 20562 11390 20562 11390 0 _0629_
rlabel metal2 21758 10642 21758 10642 0 _0630_
rlabel metal1 20102 11050 20102 11050 0 _0631_
rlabel metal1 18630 11118 18630 11118 0 _0632_
rlabel metal1 17250 10608 17250 10608 0 _0633_
rlabel metal1 17526 11084 17526 11084 0 _0634_
rlabel metal1 17250 10982 17250 10982 0 _0635_
rlabel via1 17066 10234 17066 10234 0 _0636_
rlabel metal2 17066 8772 17066 8772 0 _0637_
rlabel metal2 17618 9146 17618 9146 0 _0638_
rlabel metal2 17894 9418 17894 9418 0 _0639_
rlabel metal1 18722 10064 18722 10064 0 _0640_
rlabel metal2 18170 10370 18170 10370 0 _0641_
rlabel metal2 7038 9947 7038 9947 0 _0642_
rlabel metal1 6992 8398 6992 8398 0 _0643_
rlabel metal2 4462 7514 4462 7514 0 _0644_
rlabel metal1 6210 7854 6210 7854 0 _0645_
rlabel metal1 5996 7412 5996 7412 0 _0646_
rlabel metal2 6578 6766 6578 6766 0 _0647_
rlabel metal1 5382 7990 5382 7990 0 _0648_
rlabel metal1 6808 8058 6808 8058 0 _0649_
rlabel metal1 5474 10506 5474 10506 0 _0650_
rlabel metal1 3450 10642 3450 10642 0 _0651_
rlabel metal1 2254 11084 2254 11084 0 _0652_
rlabel metal1 3910 10778 3910 10778 0 _0653_
rlabel metal1 1610 11186 1610 11186 0 _0654_
rlabel metal1 4324 11186 4324 11186 0 _0655_
rlabel metal2 3542 13124 3542 13124 0 _0656_
rlabel metal1 4738 11322 4738 11322 0 _0657_
rlabel metal1 5428 15402 5428 15402 0 _0658_
rlabel metal1 4600 15470 4600 15470 0 _0659_
rlabel metal1 3957 17306 3957 17306 0 _0660_
rlabel metal1 4646 15606 4646 15606 0 _0661_
rlabel metal1 4830 16150 4830 16150 0 _0662_
rlabel metal2 4186 17714 4186 17714 0 _0663_
rlabel metal1 4301 17034 4301 17034 0 _0664_
rlabel metal1 3542 17612 3542 17612 0 _0665_
rlabel metal1 2254 17850 2254 17850 0 _0666_
rlabel metal1 4784 18734 4784 18734 0 _0667_
rlabel metal1 4922 17646 4922 17646 0 _0668_
rlabel metal2 5382 16932 5382 16932 0 _0669_
rlabel metal1 9154 16116 9154 16116 0 _0670_
rlabel metal2 8878 16354 8878 16354 0 _0671_
rlabel metal1 9430 17170 9430 17170 0 _0672_
rlabel metal1 10672 15538 10672 15538 0 _0673_
rlabel metal1 10212 16422 10212 16422 0 _0674_
rlabel metal2 10442 17612 10442 17612 0 _0675_
rlabel metal2 10994 16252 10994 16252 0 _0676_
rlabel metal2 11362 16320 11362 16320 0 _0677_
rlabel metal1 10810 17238 10810 17238 0 _0678_
rlabel metal2 11822 15776 11822 15776 0 _0679_
rlabel via1 20280 16082 20280 16082 0 _0680_
rlabel metal1 19182 14042 19182 14042 0 _0681_
rlabel metal1 17894 14348 17894 14348 0 _0682_
rlabel metal1 19458 14518 19458 14518 0 _0683_
rlabel metal1 18860 15946 18860 15946 0 _0684_
rlabel metal2 17342 15300 17342 15300 0 _0685_
rlabel metal1 18262 15470 18262 15470 0 _0686_
rlabel metal1 18170 14518 18170 14518 0 _0687_
rlabel metal1 18400 15674 18400 15674 0 _0688_
rlabel metal1 17848 16014 17848 16014 0 _0689_
rlabel metal1 17618 15946 17618 15946 0 _0690_
rlabel metal1 17020 15878 17020 15878 0 _0691_
rlabel metal2 20378 16286 20378 16286 0 _0692_
rlabel metal1 21505 16218 21505 16218 0 _0693_
rlabel metal1 22356 14926 22356 14926 0 _0694_
rlabel via1 21942 17170 21942 17170 0 _0695_
rlabel viali 21942 17646 21942 17646 0 _0696_
rlabel metal2 22126 16796 22126 16796 0 _0697_
rlabel metal2 22402 16796 22402 16796 0 _0698_
rlabel metal2 21942 18054 21942 18054 0 _0699_
rlabel metal1 22586 18190 22586 18190 0 _0700_
rlabel metal2 21666 18462 21666 18462 0 _0701_
rlabel metal1 23092 15402 23092 15402 0 _0702_
rlabel metal2 18170 16932 18170 16932 0 _0703_
rlabel metal2 17986 15028 17986 15028 0 _0704_
rlabel metal2 17434 14042 17434 14042 0 _0705_
rlabel via2 18630 14467 18630 14467 0 _0706_
rlabel metal1 20148 14042 20148 14042 0 _0707_
rlabel metal1 16514 14042 16514 14042 0 _0708_
rlabel metal1 18998 17306 18998 17306 0 _0709_
rlabel metal2 15962 15334 15962 15334 0 _0710_
rlabel metal2 8970 15844 8970 15844 0 _0711_
rlabel metal1 9982 16048 9982 16048 0 _0712_
rlabel metal2 10534 15844 10534 15844 0 _0713_
rlabel metal2 10258 16694 10258 16694 0 _0714_
rlabel metal1 12558 17136 12558 17136 0 _0715_
rlabel metal1 9660 17102 9660 17102 0 _0716_
rlabel metal1 8786 17170 8786 17170 0 _0717_
rlabel metal2 12926 16796 12926 16796 0 _0718_
rlabel metal2 12742 16762 12742 16762 0 _0719_
rlabel metal1 11546 16218 11546 16218 0 _0720_
rlabel metal1 7728 15470 7728 15470 0 _0721_
rlabel metal2 3358 17918 3358 17918 0 _0722_
rlabel metal1 3726 17714 3726 17714 0 _0723_
rlabel metal1 4462 18258 4462 18258 0 _0724_
rlabel metal2 4278 18462 4278 18462 0 _0725_
rlabel metal2 5106 19108 5106 19108 0 _0726_
rlabel metal1 3956 17850 3956 17850 0 _0727_
rlabel metal1 2576 18394 2576 18394 0 _0728_
rlabel metal1 3634 15504 3634 15504 0 _0729_
rlabel metal2 3634 15844 3634 15844 0 _0730_
rlabel metal2 4922 10234 4922 10234 0 _0731_
rlabel metal1 4094 10234 4094 10234 0 _0732_
rlabel metal2 2714 10914 2714 10914 0 _0733_
rlabel metal1 2024 11186 2024 11186 0 _0734_
rlabel metal1 2576 11322 2576 11322 0 _0735_
rlabel metal1 3634 13226 3634 13226 0 _0736_
rlabel metal1 2070 11322 2070 11322 0 _0737_
rlabel metal2 2714 9146 2714 9146 0 _0738_
rlabel metal1 5290 10030 5290 10030 0 _0739_
rlabel metal1 4876 9690 4876 9690 0 _0740_
rlabel metal1 6164 7310 6164 7310 0 _0741_
rlabel metal1 4784 7446 4784 7446 0 _0742_
rlabel metal1 4646 7344 4646 7344 0 _0743_
rlabel metal1 4600 6834 4600 6834 0 _0744_
rlabel metal1 4968 5338 4968 5338 0 _0745_
rlabel metal1 3128 7514 3128 7514 0 _0746_
rlabel metal2 7038 5916 7038 5916 0 _0747_
rlabel metal1 7084 8466 7084 8466 0 _0748_
rlabel metal1 17342 11152 17342 11152 0 _0749_
rlabel metal2 17434 10812 17434 10812 0 _0750_
rlabel metal2 17434 9690 17434 9690 0 _0751_
rlabel metal2 16974 9316 16974 9316 0 _0752_
rlabel metal2 15594 9146 15594 9146 0 _0753_
rlabel metal1 18768 8602 18768 8602 0 _0754_
rlabel metal2 17526 11968 17526 11968 0 _0755_
rlabel metal1 19734 11254 19734 11254 0 _0756_
rlabel metal1 19642 11322 19642 11322 0 _0757_
rlabel metal1 21528 9690 21528 9690 0 _0758_
rlabel metal1 22678 9962 22678 9962 0 _0759_
rlabel metal1 21068 11662 21068 11662 0 _0760_
rlabel metal1 24196 12138 24196 12138 0 _0761_
rlabel metal1 28198 10608 28198 10608 0 _0762_
rlabel metal1 27692 12750 27692 12750 0 _0763_
rlabel metal1 26404 12750 26404 12750 0 _0764_
rlabel metal2 27186 13668 27186 13668 0 _0765_
rlabel metal1 28014 15334 28014 15334 0 _0766_
rlabel metal1 26496 14926 26496 14926 0 _0767_
rlabel metal2 25070 17306 25070 17306 0 _0768_
rlabel metal1 26956 17578 26956 17578 0 _0769_
rlabel metal2 27738 19924 27738 19924 0 _0770_
rlabel metal1 26312 19278 26312 19278 0 _0771_
rlabel metal1 25484 21658 25484 21658 0 _0772_
rlabel metal2 27002 21801 27002 21801 0 _0773_
rlabel metal2 27738 23460 27738 23460 0 _0774_
rlabel metal1 26956 24582 26956 24582 0 _0775_
rlabel metal1 27416 25466 27416 25466 0 _0776_
rlabel metal1 25652 27370 25652 27370 0 _0777_
rlabel metal1 25162 27370 25162 27370 0 _0778_
rlabel metal1 23744 26282 23744 26282 0 _0779_
rlabel metal1 23736 25262 23736 25262 0 _0780_
rlabel metal2 16238 26146 16238 26146 0 _0781_
rlabel metal1 16514 25262 16514 25262 0 _0782_
rlabel metal2 15870 25568 15870 25568 0 _0783_
rlabel metal1 15318 25330 15318 25330 0 _0784_
rlabel metal1 16652 25466 16652 25466 0 _0785_
rlabel metal2 16882 25398 16882 25398 0 _0786_
rlabel metal1 17434 26316 17434 26316 0 _0787_
rlabel metal1 16330 26384 16330 26384 0 _0788_
rlabel metal1 16054 26248 16054 26248 0 _0789_
rlabel metal1 15962 26350 15962 26350 0 _0790_
rlabel metal1 15732 26350 15732 26350 0 _0791_
rlabel metal2 13110 25602 13110 25602 0 _0792_
rlabel metal2 13386 25670 13386 25670 0 _0793_
rlabel metal1 13616 26010 13616 26010 0 _0794_
rlabel metal1 10948 26350 10948 26350 0 _0795_
rlabel metal1 11822 25398 11822 25398 0 _0796_
rlabel metal1 9614 25908 9614 25908 0 _0797_
rlabel metal2 9890 26044 9890 26044 0 _0798_
rlabel metal2 9982 25568 9982 25568 0 _0799_
rlabel metal1 12834 25840 12834 25840 0 _0800_
rlabel metal2 10994 26044 10994 26044 0 _0801_
rlabel metal1 10580 26010 10580 26010 0 _0802_
rlabel metal2 12650 26656 12650 26656 0 _0803_
rlabel metal1 13294 25840 13294 25840 0 _0804_
rlabel metal1 18814 5168 18814 5168 0 _0805_
rlabel metal2 22494 4964 22494 4964 0 _0806_
rlabel metal1 22816 4726 22816 4726 0 _0807_
rlabel metal1 22586 4794 22586 4794 0 _0808_
rlabel metal1 21298 5338 21298 5338 0 _0809_
rlabel metal1 20746 5202 20746 5202 0 _0810_
rlabel metal2 20102 5372 20102 5372 0 _0811_
rlabel metal1 18906 5236 18906 5236 0 _0812_
rlabel metal2 18630 5542 18630 5542 0 _0813_
rlabel metal2 16514 5610 16514 5610 0 _0814_
rlabel metal2 16882 5508 16882 5508 0 _0815_
rlabel metal1 15042 5882 15042 5882 0 _0816_
rlabel metal2 12650 6596 12650 6596 0 _0817_
rlabel metal1 13708 5882 13708 5882 0 _0818_
rlabel metal2 14122 6460 14122 6460 0 _0819_
rlabel metal1 13156 6426 13156 6426 0 _0820_
rlabel metal1 13202 6732 13202 6732 0 _0821_
rlabel metal1 12788 6970 12788 6970 0 _0822_
rlabel metal2 12650 9044 12650 9044 0 _0823_
rlabel metal1 12558 7514 12558 7514 0 _0824_
rlabel metal2 14030 14178 14030 14178 0 _0825_
rlabel metal2 13478 13770 13478 13770 0 _0826_
rlabel metal1 13570 13906 13570 13906 0 _0827_
rlabel metal1 13064 13294 13064 13294 0 _0828_
rlabel metal2 12926 12682 12926 12682 0 _0829_
rlabel metal2 12834 10948 12834 10948 0 _0830_
rlabel metal2 13018 11968 13018 11968 0 _0831_
rlabel metal2 12558 11322 12558 11322 0 _0832_
rlabel metal2 13110 11900 13110 11900 0 _0833_
rlabel metal1 13432 12206 13432 12206 0 _0834_
rlabel metal2 12650 17204 12650 17204 0 _0835_
rlabel metal2 11914 25670 11914 25670 0 _0836_
rlabel metal1 12006 25704 12006 25704 0 _0837_
rlabel metal2 12466 26112 12466 26112 0 _0838_
rlabel metal1 12558 25704 12558 25704 0 _0839_
rlabel metal2 12650 25721 12650 25721 0 _0840_
rlabel metal2 17618 25636 17618 25636 0 _0841_
rlabel metal2 15962 26486 15962 26486 0 _0842_
rlabel metal1 15778 25908 15778 25908 0 _0843_
rlabel metal2 15226 26384 15226 26384 0 _0844_
rlabel metal1 14628 26010 14628 26010 0 _0845_
rlabel metal2 15318 26554 15318 26554 0 _0846_
rlabel metal1 23184 2346 23184 2346 0 _0847_
rlabel metal1 23368 2618 23368 2618 0 _0848_
rlabel via1 23422 2346 23422 2346 0 _0849_
rlabel metal1 21896 3094 21896 3094 0 _0850_
rlabel metal1 20792 3434 20792 3434 0 _0851_
rlabel metal1 19412 3570 19412 3570 0 _0852_
rlabel metal1 20056 3706 20056 3706 0 _0853_
rlabel metal2 18078 3808 18078 3808 0 _0854_
rlabel metal1 18684 3366 18684 3366 0 _0855_
rlabel metal1 16468 3638 16468 3638 0 _0856_
rlabel metal2 16606 3808 16606 3808 0 _0857_
rlabel metal1 14720 4046 14720 4046 0 _0858_
rlabel metal1 15640 3094 15640 3094 0 _0859_
rlabel metal1 12006 4114 12006 4114 0 _0860_
rlabel metal1 13508 3434 13508 3434 0 _0861_
rlabel metal1 11040 4182 11040 4182 0 _0862_
rlabel metal1 10902 3706 10902 3706 0 _0863_
rlabel metal1 13340 10642 13340 10642 0 _0864_
rlabel metal1 11730 3944 11730 3944 0 _0865_
rlabel metal1 14122 11696 14122 11696 0 _0866_
rlabel metal1 13624 9894 13624 9894 0 _0867_
rlabel metal2 14214 11934 14214 11934 0 _0868_
rlabel metal1 14582 11560 14582 11560 0 _0869_
rlabel metal2 13386 11169 13386 11169 0 _0870_
rlabel metal1 14812 12342 14812 12342 0 _0871_
rlabel metal1 6946 15028 6946 15028 0 _0872_
rlabel viali 6179 12172 6179 12172 0 _0873_
rlabel metal1 6670 14518 6670 14518 0 _0874_
rlabel metal2 6762 14688 6762 14688 0 _0875_
rlabel metal1 4876 13906 4876 13906 0 _0876_
rlabel metal1 5060 13702 5060 13702 0 _0877_
rlabel metal2 4186 23970 4186 23970 0 _0878_
rlabel metal1 4592 21862 4592 21862 0 _0879_
rlabel metal1 4692 24310 4692 24310 0 _0880_
rlabel metal1 4600 24378 4600 24378 0 _0881_
rlabel metal2 4738 24378 4738 24378 0 _0882_
rlabel metal1 4508 25466 4508 25466 0 _0883_
rlabel via1 6854 27438 6854 27438 0 _0884_
rlabel metal1 6616 27098 6616 27098 0 _0885_
rlabel metal2 7590 27812 7590 27812 0 _0886_
rlabel metal1 7820 27642 7820 27642 0 _0887_
rlabel metal1 13570 27472 13570 27472 0 _0888_
rlabel metal1 7498 28594 7498 28594 0 _0889_
rlabel metal2 10074 27846 10074 27846 0 _0890_
rlabel metal2 12742 28356 12742 28356 0 _0891_
rlabel metal1 10948 27642 10948 27642 0 _0892_
rlabel metal1 14674 27438 14674 27438 0 _0893_
rlabel metal1 14122 27438 14122 27438 0 _0894_
rlabel metal1 14812 27642 14812 27642 0 _0895_
rlabel metal1 14674 27914 14674 27914 0 _0896_
rlabel metal1 16008 27642 16008 27642 0 _0897_
rlabel metal1 17572 28526 17572 28526 0 _0898_
rlabel metal1 17940 27370 17940 27370 0 _0899_
rlabel metal1 17572 27574 17572 27574 0 _0900_
rlabel metal1 19688 27846 19688 27846 0 _0901_
rlabel metal1 19466 28186 19466 28186 0 _0902_
rlabel metal1 19688 27302 19688 27302 0 _0903_
rlabel metal1 19320 27574 19320 27574 0 _0904_
rlabel metal1 20424 26554 20424 26554 0 _0905_
rlabel metal1 20202 26214 20202 26214 0 _0906_
rlabel metal1 24150 20774 24150 20774 0 _0907_
rlabel metal2 23138 21182 23138 21182 0 _0908_
rlabel metal1 12880 24038 12880 24038 0 _0909_
rlabel metal1 10626 23086 10626 23086 0 _0910_
rlabel metal1 7958 23562 7958 23562 0 _0911_
rlabel metal1 12558 23052 12558 23052 0 _0912_
rlabel metal2 11178 23426 11178 23426 0 _0913_
rlabel metal2 10810 23868 10810 23868 0 _0914_
rlabel metal1 11454 23698 11454 23698 0 _0915_
rlabel metal1 10258 23766 10258 23766 0 _0916_
rlabel metal1 11730 23664 11730 23664 0 _0917_
rlabel metal1 12604 23698 12604 23698 0 _0918_
rlabel metal1 14122 23800 14122 23800 0 _0919_
rlabel metal1 21482 6358 21482 6358 0 _0920_
rlabel metal2 24794 5882 24794 5882 0 _0921_
rlabel metal2 24978 5882 24978 5882 0 _0922_
rlabel metal2 21482 5950 21482 5950 0 _0923_
rlabel metal1 21344 5814 21344 5814 0 _0924_
rlabel metal1 19182 5338 19182 5338 0 _0925_
rlabel metal2 18538 4998 18538 4998 0 _0926_
rlabel metal1 17848 5202 17848 5202 0 _0927_
rlabel metal1 16192 5270 16192 5270 0 _0928_
rlabel metal2 14858 4998 14858 4998 0 _0929_
rlabel metal1 14122 4794 14122 4794 0 _0930_
rlabel metal1 13386 5236 13386 5236 0 _0931_
rlabel metal2 14168 5338 14168 5338 0 _0932_
rlabel metal1 13708 7378 13708 7378 0 _0933_
rlabel metal1 14444 7514 14444 7514 0 _0934_
rlabel metal1 13892 8602 13892 8602 0 _0935_
rlabel metal1 12006 13294 12006 13294 0 _0936_
rlabel metal2 10626 13770 10626 13770 0 _0937_
rlabel metal1 10626 13872 10626 13872 0 _0938_
rlabel metal1 11500 13498 11500 13498 0 _0939_
rlabel metal1 10534 13328 10534 13328 0 _0940_
rlabel metal1 11454 13294 11454 13294 0 _0941_
rlabel metal1 15364 15402 15364 15402 0 clk
rlabel metal1 16606 15674 16606 15674 0 clknet_0_clk
rlabel metal1 2208 13838 2208 13838 0 clknet_3_0__leaf_clk
rlabel metal1 14674 13362 14674 13362 0 clknet_3_1__leaf_clk
rlabel metal1 1702 16150 1702 16150 0 clknet_3_2__leaf_clk
rlabel metal2 12650 28560 12650 28560 0 clknet_3_3__leaf_clk
rlabel metal2 20654 13124 20654 13124 0 clknet_3_4__leaf_clk
rlabel metal2 27646 13838 27646 13838 0 clknet_3_5__leaf_clk
rlabel metal1 21344 22066 21344 22066 0 clknet_3_6__leaf_clk
rlabel metal2 27600 21522 27600 21522 0 clknet_3_7__leaf_clk
rlabel metal1 24104 4590 24104 4590 0 fast_pwm_inst.pwm_counter\[0\]
rlabel metal1 13294 7854 13294 7854 0 fast_pwm_inst.pwm_counter\[10\]
rlabel metal1 14536 10642 14536 10642 0 fast_pwm_inst.pwm_counter\[11\]
rlabel metal2 9062 11900 9062 11900 0 fast_pwm_inst.pwm_counter\[12\]
rlabel metal1 8786 12784 8786 12784 0 fast_pwm_inst.pwm_counter\[13\]
rlabel metal1 10810 13260 10810 13260 0 fast_pwm_inst.pwm_counter\[14\]
rlabel metal1 13524 14382 13524 14382 0 fast_pwm_inst.pwm_counter\[15\]
rlabel via1 7498 23086 7498 23086 0 fast_pwm_inst.pwm_counter\[16\]
rlabel metal1 5658 22984 5658 22984 0 fast_pwm_inst.pwm_counter\[17\]
rlabel metal1 5428 26010 5428 26010 0 fast_pwm_inst.pwm_counter\[18\]
rlabel metal1 7314 23664 7314 23664 0 fast_pwm_inst.pwm_counter\[19\]
rlabel metal2 23782 3332 23782 3332 0 fast_pwm_inst.pwm_counter\[1\]
rlabel metal1 9729 26962 9729 26962 0 fast_pwm_inst.pwm_counter\[20\]
rlabel via1 7498 27914 7498 27914 0 fast_pwm_inst.pwm_counter\[21\]
rlabel metal2 13294 24684 13294 24684 0 fast_pwm_inst.pwm_counter\[22\]
rlabel metal1 13018 25262 13018 25262 0 fast_pwm_inst.pwm_counter\[23\]
rlabel metal2 13202 28050 13202 28050 0 fast_pwm_inst.pwm_counter\[24\]
rlabel metal2 15502 28458 15502 28458 0 fast_pwm_inst.pwm_counter\[25\]
rlabel metal1 15502 27370 15502 27370 0 fast_pwm_inst.pwm_counter\[26\]
rlabel metal1 18722 29274 18722 29274 0 fast_pwm_inst.pwm_counter\[27\]
rlabel metal1 21482 24106 21482 24106 0 fast_pwm_inst.pwm_counter\[28\]
rlabel metal1 19826 24820 19826 24820 0 fast_pwm_inst.pwm_counter\[29\]
rlabel metal1 21114 5168 21114 5168 0 fast_pwm_inst.pwm_counter\[2\]
rlabel metal1 20378 26350 20378 26350 0 fast_pwm_inst.pwm_counter\[30\]
rlabel metal1 19274 25942 19274 25942 0 fast_pwm_inst.pwm_counter\[31\]
rlabel metal1 21160 3910 21160 3910 0 fast_pwm_inst.pwm_counter\[3\]
rlabel metal1 18032 4114 18032 4114 0 fast_pwm_inst.pwm_counter\[4\]
rlabel metal2 17618 3162 17618 3162 0 fast_pwm_inst.pwm_counter\[5\]
rlabel metal2 16146 3230 16146 3230 0 fast_pwm_inst.pwm_counter\[6\]
rlabel metal1 14950 4114 14950 4114 0 fast_pwm_inst.pwm_counter\[7\]
rlabel metal1 13018 6868 13018 6868 0 fast_pwm_inst.pwm_counter\[8\]
rlabel metal1 12282 4590 12282 4590 0 fast_pwm_inst.pwm_counter\[9\]
rlabel metal2 22954 21692 22954 21692 0 fast_pwm_inst.pwm_outa
rlabel metal1 24012 22406 24012 22406 0 fast_pwm_inst.pwm_outb
rlabel metal2 25438 22882 25438 22882 0 irq_timer_normal
rlabel metal1 14674 8840 14674 8840 0 net1
rlabel via2 1702 10659 1702 10659 0 net10
rlabel metal1 1886 3060 1886 3060 0 net100
rlabel metal1 24932 20774 24932 20774 0 net101
rlabel metal1 28244 16558 28244 16558 0 net102
rlabel metal1 20654 26520 20654 26520 0 net11
rlabel metal1 2024 24582 2024 24582 0 net12
rlabel metal1 2231 18802 2231 18802 0 net13
rlabel metal1 7774 18734 7774 18734 0 net14
rlabel metal2 1610 16082 1610 16082 0 net15
rlabel metal1 14168 24106 14168 24106 0 net16
rlabel metal1 14582 21998 14582 21998 0 net17
rlabel via1 15136 19822 15136 19822 0 net18
rlabel metal1 19458 21930 19458 21930 0 net19
rlabel metal1 1748 21386 1748 21386 0 net2
rlabel metal1 23529 2278 23529 2278 0 net20
rlabel metal2 21482 17867 21482 17867 0 net21
rlabel metal1 21390 20298 21390 20298 0 net22
rlabel metal2 23874 8602 23874 8602 0 net23
rlabel metal1 21206 19856 21206 19856 0 net24
rlabel via2 1702 19805 1702 19805 0 net25
rlabel metal2 22310 17238 22310 17238 0 net26
rlabel metal2 13294 2142 13294 2142 0 net27
rlabel metal2 18538 7055 18538 7055 0 net28
rlabel metal2 17618 7463 17618 7463 0 net29
rlabel metal2 27278 2040 27278 2040 0 net3
rlabel metal1 8556 2414 8556 2414 0 net30
rlabel metal1 5474 2380 5474 2380 0 net31
rlabel metal1 2231 6222 2231 6222 0 net32
rlabel metal1 27278 7786 27278 7786 0 net33
rlabel metal2 13754 7905 13754 7905 0 net34
rlabel metal2 29210 1972 29210 1972 0 net35
rlabel metal2 23690 2550 23690 2550 0 net36
rlabel metal1 26174 14518 26174 14518 0 net37
rlabel metal2 21942 11424 21942 11424 0 net38
rlabel metal2 12006 21726 12006 21726 0 net39
rlabel metal2 15732 25364 15732 25364 0 net4
rlabel metal1 11730 30022 11730 30022 0 net40
rlabel metal1 20010 24650 20010 24650 0 net41
rlabel metal2 1610 4862 1610 4862 0 net42
rlabel metal1 8510 2618 8510 2618 0 net43
rlabel metal1 24610 7888 24610 7888 0 net44
rlabel via1 9248 20434 9248 20434 0 net45
rlabel metal1 16882 30158 16882 30158 0 net46
rlabel metal1 2231 23630 2231 23630 0 net47
rlabel metal1 9522 30158 9522 30158 0 net48
rlabel via2 14214 21981 14214 21981 0 net49
rlabel metal1 1840 30158 1840 30158 0 net5
rlabel metal1 14858 21998 14858 21998 0 net50
rlabel metal2 16882 21471 16882 21471 0 net51
rlabel metal1 17020 21998 17020 21998 0 net52
rlabel metal1 12006 2618 12006 2618 0 net53
rlabel metal1 18630 18666 18630 18666 0 net54
rlabel metal1 29532 20774 29532 20774 0 net55
rlabel metal1 18676 18938 18676 18938 0 net56
rlabel metal1 18308 20434 18308 20434 0 net57
rlabel metal1 20194 7378 20194 7378 0 net58
rlabel metal1 18722 4522 18722 4522 0 net59
rlabel metal1 16422 12682 16422 12682 0 net6
rlabel metal2 1610 3094 1610 3094 0 net60
rlabel metal1 18906 2550 18906 2550 0 net61
rlabel metal1 2346 2550 2346 2550 0 net62
rlabel metal2 10442 4148 10442 4148 0 net63
rlabel metal2 28198 2142 28198 2142 0 net64
rlabel metal1 23000 2618 23000 2618 0 net65
rlabel metal1 1886 26282 1886 26282 0 net66
rlabel metal1 19550 3570 19550 3570 0 net67
rlabel metal1 12742 10982 12742 10982 0 net68
rlabel via1 13385 13906 13385 13906 0 net69
rlabel metal1 5014 2278 5014 2278 0 net7
rlabel metal1 20470 13906 20470 13906 0 net70
rlabel via2 25898 2397 25898 2397 0 net71
rlabel metal2 13938 21148 13938 21148 0 net72
rlabel metal1 14260 2618 14260 2618 0 net73
rlabel metal1 9568 20366 9568 20366 0 net74
rlabel metal1 2530 13804 2530 13804 0 net75
rlabel metal2 1610 2108 1610 2108 0 net76
rlabel via2 18906 2261 18906 2261 0 net77
rlabel metal1 10994 22644 10994 22644 0 net78
rlabel metal2 13570 29818 13570 29818 0 net79
rlabel metal2 15962 24990 15962 24990 0 net8
rlabel metal2 12834 20145 12834 20145 0 net80
rlabel metal1 14490 19380 14490 19380 0 net81
rlabel via2 5014 2533 5014 2533 0 net82
rlabel metal1 1840 18258 1840 18258 0 net83
rlabel metal2 27922 24905 27922 24905 0 net84
rlabel metal1 18078 18768 18078 18768 0 net85
rlabel metal1 15870 2380 15870 2380 0 net86
rlabel metal2 28152 12420 28152 12420 0 net87
rlabel metal1 18998 4998 18998 4998 0 net88
rlabel metal2 18354 18326 18354 18326 0 net89
rlabel via2 6394 22627 6394 22627 0 net9
rlabel metal2 1978 8959 1978 8959 0 net90
rlabel metal1 18584 2618 18584 2618 0 net91
rlabel metal1 13156 2278 13156 2278 0 net92
rlabel metal2 16238 5984 16238 5984 0 net93
rlabel metal1 19918 5814 19918 5814 0 net94
rlabel metal1 14490 5610 14490 5610 0 net95
rlabel metal1 13570 6324 13570 6324 0 net96
rlabel metal2 23966 21529 23966 21529 0 net97
rlabel metal2 2714 26554 2714 26554 0 net98
rlabel metal1 2300 13294 2300 13294 0 net99
rlabel metal1 26128 11118 26128 11118 0 normal_mode_inst.timer_cnt\[0\]
rlabel metal2 25622 16966 25622 16966 0 normal_mode_inst.timer_cnt\[10\]
rlabel metal1 26312 17170 26312 17170 0 normal_mode_inst.timer_cnt\[11\]
rlabel metal1 27876 17306 27876 17306 0 normal_mode_inst.timer_cnt\[12\]
rlabel metal2 27554 18530 27554 18530 0 normal_mode_inst.timer_cnt\[13\]
rlabel metal2 27554 20230 27554 20230 0 normal_mode_inst.timer_cnt\[14\]
rlabel metal1 27278 19958 27278 19958 0 normal_mode_inst.timer_cnt\[15\]
rlabel metal1 26404 21522 26404 21522 0 normal_mode_inst.timer_cnt\[16\]
rlabel metal1 25714 21862 25714 21862 0 normal_mode_inst.timer_cnt\[17\]
rlabel metal2 27186 21760 27186 21760 0 normal_mode_inst.timer_cnt\[18\]
rlabel metal1 27692 23018 27692 23018 0 normal_mode_inst.timer_cnt\[19\]
rlabel metal2 27738 9962 27738 9962 0 normal_mode_inst.timer_cnt\[1\]
rlabel metal1 27692 23698 27692 23698 0 normal_mode_inst.timer_cnt\[20\]
rlabel metal1 27324 24378 27324 24378 0 normal_mode_inst.timer_cnt\[21\]
rlabel metal1 27370 25976 27370 25976 0 normal_mode_inst.timer_cnt\[22\]
rlabel metal2 28014 26894 28014 26894 0 normal_mode_inst.timer_cnt\[23\]
rlabel metal1 27002 26418 27002 26418 0 normal_mode_inst.timer_cnt\[24\]
rlabel metal2 27186 28220 27186 28220 0 normal_mode_inst.timer_cnt\[25\]
rlabel metal2 25806 28050 25806 28050 0 normal_mode_inst.timer_cnt\[26\]
rlabel metal2 24242 28220 24242 28220 0 normal_mode_inst.timer_cnt\[27\]
rlabel metal2 23506 27778 23506 27778 0 normal_mode_inst.timer_cnt\[28\]
rlabel metal2 23506 26520 23506 26520 0 normal_mode_inst.timer_cnt\[29\]
rlabel metal1 27554 9928 27554 9928 0 normal_mode_inst.timer_cnt\[2\]
rlabel metal2 24058 24990 24058 24990 0 normal_mode_inst.timer_cnt\[30\]
rlabel metal2 23598 24990 23598 24990 0 normal_mode_inst.timer_cnt\[31\]
rlabel metal2 28290 11322 28290 11322 0 normal_mode_inst.timer_cnt\[3\]
rlabel metal1 27370 12818 27370 12818 0 normal_mode_inst.timer_cnt\[4\]
rlabel metal2 27186 12886 27186 12886 0 normal_mode_inst.timer_cnt\[5\]
rlabel metal1 27416 13294 27416 13294 0 normal_mode_inst.timer_cnt\[6\]
rlabel metal1 28980 14858 28980 14858 0 normal_mode_inst.timer_cnt\[7\]
rlabel metal1 27416 16082 27416 16082 0 normal_mode_inst.timer_cnt\[8\]
rlabel metal2 27462 14756 27462 14756 0 normal_mode_inst.timer_cnt\[9\]
rlabel metal1 22126 13872 22126 13872 0 phase_pwm_inst.counter\[0\]
rlabel metal1 8050 7412 8050 7412 0 phase_pwm_inst.counter\[10\]
rlabel metal2 5934 5406 5934 5406 0 phase_pwm_inst.counter\[11\]
rlabel metal2 10626 10302 10626 10302 0 phase_pwm_inst.counter\[12\]
rlabel metal2 2622 10931 2622 10931 0 phase_pwm_inst.counter\[13\]
rlabel metal1 7820 13158 7820 13158 0 phase_pwm_inst.counter\[14\]
rlabel metal2 7222 13328 7222 13328 0 phase_pwm_inst.counter\[15\]
rlabel metal1 9982 19992 9982 19992 0 phase_pwm_inst.counter\[16\]
rlabel metal2 7682 22372 7682 22372 0 phase_pwm_inst.counter\[17\]
rlabel metal1 5750 17646 5750 17646 0 phase_pwm_inst.counter\[18\]
rlabel metal1 8970 19856 8970 19856 0 phase_pwm_inst.counter\[19\]
rlabel metal2 21850 7684 21850 7684 0 phase_pwm_inst.counter\[1\]
rlabel metal1 9384 21998 9384 21998 0 phase_pwm_inst.counter\[20\]
rlabel metal1 10810 18360 10810 18360 0 phase_pwm_inst.counter\[21\]
rlabel metal1 13938 17170 13938 17170 0 phase_pwm_inst.counter\[22\]
rlabel metal1 13110 21488 13110 21488 0 phase_pwm_inst.counter\[23\]
rlabel metal1 14582 19890 14582 19890 0 phase_pwm_inst.counter\[24\]
rlabel metal1 14950 21488 14950 21488 0 phase_pwm_inst.counter\[25\]
rlabel metal2 19090 21250 19090 21250 0 phase_pwm_inst.counter\[26\]
rlabel metal1 17388 19346 17388 19346 0 phase_pwm_inst.counter\[27\]
rlabel metal2 21942 19890 21942 19890 0 phase_pwm_inst.counter\[28\]
rlabel metal2 21850 18666 21850 18666 0 phase_pwm_inst.counter\[29\]
rlabel metal1 21666 7752 21666 7752 0 phase_pwm_inst.counter\[2\]
rlabel metal1 22862 18326 22862 18326 0 phase_pwm_inst.counter\[30\]
rlabel metal1 21482 16626 21482 16626 0 phase_pwm_inst.counter\[31\]
rlabel metal1 20608 9554 20608 9554 0 phase_pwm_inst.counter\[3\]
rlabel metal1 20056 12206 20056 12206 0 phase_pwm_inst.counter\[4\]
rlabel metal1 18170 12954 18170 12954 0 phase_pwm_inst.counter\[5\]
rlabel metal2 19274 9588 19274 9588 0 phase_pwm_inst.counter\[6\]
rlabel metal1 17158 10030 17158 10030 0 phase_pwm_inst.counter\[7\]
rlabel metal2 13018 9180 13018 9180 0 phase_pwm_inst.counter\[8\]
rlabel metal2 8050 5508 8050 5508 0 phase_pwm_inst.counter\[9\]
rlabel metal1 20470 13294 20470 13294 0 phase_pwm_inst.direction
rlabel metal2 23230 21318 23230 21318 0 phase_pwm_inst.pwm_outa
rlabel metal2 24518 20740 24518 20740 0 phase_pwm_inst.pwm_outb
rlabel metal3 1050 28628 1050 28628 0 reset
rlabel via2 28474 16405 28474 16405 0 timer_interrupt
<< properties >>
string FIXED_BBOX 0 0 30903 33047
<< end >>
