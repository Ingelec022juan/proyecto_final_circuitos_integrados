* NGSPICE file created from Timer_PWM_Generator.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt Timer_PWM_Generator PWM_CNTA[0] PWM_CNTA[10] PWM_CNTA[11] PWM_CNTA[12] PWM_CNTA[13]
+ PWM_CNTA[14] PWM_CNTA[15] PWM_CNTA[16] PWM_CNTA[17] PWM_CNTA[18] PWM_CNTA[19] PWM_CNTA[1]
+ PWM_CNTA[20] PWM_CNTA[21] PWM_CNTA[22] PWM_CNTA[23] PWM_CNTA[24] PWM_CNTA[25] PWM_CNTA[26]
+ PWM_CNTA[27] PWM_CNTA[28] PWM_CNTA[29] PWM_CNTA[2] PWM_CNTA[30] PWM_CNTA[31] PWM_CNTA[3]
+ PWM_CNTA[4] PWM_CNTA[5] PWM_CNTA[6] PWM_CNTA[7] PWM_CNTA[8] PWM_CNTA[9] PWM_CNTB[0]
+ PWM_CNTB[10] PWM_CNTB[11] PWM_CNTB[12] PWM_CNTB[13] PWM_CNTB[14] PWM_CNTB[15] PWM_CNTB[16]
+ PWM_CNTB[17] PWM_CNTB[18] PWM_CNTB[19] PWM_CNTB[1] PWM_CNTB[20] PWM_CNTB[21] PWM_CNTB[22]
+ PWM_CNTB[23] PWM_CNTB[24] PWM_CNTB[25] PWM_CNTB[26] PWM_CNTB[27] PWM_CNTB[28] PWM_CNTB[29]
+ PWM_CNTB[2] PWM_CNTB[30] PWM_CNTB[31] PWM_CNTB[3] PWM_CNTB[4] PWM_CNTB[5] PWM_CNTB[6]
+ PWM_CNTB[7] PWM_CNTB[8] PWM_CNTB[9] PWM_OUTA PWM_OUTB TIMER_TOP[0] TIMER_TOP[10]
+ TIMER_TOP[11] TIMER_TOP[12] TIMER_TOP[13] TIMER_TOP[14] TIMER_TOP[15] TIMER_TOP[16]
+ TIMER_TOP[17] TIMER_TOP[18] TIMER_TOP[19] TIMER_TOP[1] TIMER_TOP[20] TIMER_TOP[21]
+ TIMER_TOP[22] TIMER_TOP[23] TIMER_TOP[24] TIMER_TOP[25] TIMER_TOP[26] TIMER_TOP[27]
+ TIMER_TOP[28] TIMER_TOP[29] TIMER_TOP[2] TIMER_TOP[30] TIMER_TOP[31] TIMER_TOP[3]
+ TIMER_TOP[4] TIMER_TOP[5] TIMER_TOP[6] TIMER_TOP[7] TIMER_TOP[8] TIMER_TOP[9] TMR_MODE[0]
+ TMR_MODE[1] TMR_SRC[0] TMR_SRC[1] VGND VPWR clk reset timer_interrupt
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1270_ _0612_ _0650_ _0655_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__o21a_1
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1606_ _0477_ net18 VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_14_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0985_ net71 VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__inv_2
X_1468_ fast_pwm_inst.pwm_counter\[22\] _0888_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nand2_1
X_1399_ net85 _0474_ _0786_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__a21o_1
X_1537_ _0937_ _0205_ _0206_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__and4b_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1322_ normal_mode_inst.timer_cnt\[7\] normal_mode_inst.timer_cnt\[9\] normal_mode_inst.timer_cnt\[8\]
+ _0765_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__and4_1
X_1253_ _0676_ _0713_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_20_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1184_ _0659_ _0660_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__nand2_1
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0968_ phase_pwm_inst.counter\[4\] VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1871_ net99 VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
X_1940_ clknet_3_7__leaf_clk _0050_ _0123_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_14_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1305_ _0755_ phase_pwm_inst.counter\[5\] _0616_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
X_1236_ _0683_ _0705_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__xnor2_1
XFILLER_44_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1167_ phase_pwm_inst.counter\[10\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0644_ sky130_fd_sc_hd__xor2_1
X_1098_ _0571_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__and2_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1021_ fast_pwm_inst.pwm_counter\[2\] VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__inv_2
X_1785_ net97 net98 irq_timer_normal VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__nor3b_1
X_1854_ net99 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__inv_2
X_1923_ clknet_3_5__leaf_clk _0063_ _0106_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1219_ _0424_ phase_pwm_inst.direction _0680_ _0692_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_51_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1570_ _0496_ net28 net27 _0497_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__o22a_1
X_1004_ fast_pwm_inst.pwm_counter\[20\] VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__inv_2
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1768_ _0775_ _0414_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and2b_1
X_1837_ net99 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__inv_2
X_1906_ clknet_3_2__leaf_clk _0191_ _0089_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[19\]
+ sky130_fd_sc_hd__dfrtp_4
X_1699_ _0447_ net27 _0362_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__a22o_1
XFILLER_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _0288_ _0289_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__a21o_1
X_1484_ _0900_ _0847_ _0899_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__and3b_1
X_1553_ fast_pwm_inst.pwm_counter\[25\] _0503_ _0216_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ net72 VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__inv_2
X_1605_ net16 _0479_ fast_pwm_inst.pwm_counter\[24\] _0525_ VGND VGND VPWR VPWR _0275_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_8_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1536_ _0487_ net38 _0938_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__or3_1
X_1467_ fast_pwm_inst.pwm_counter\[21\] _0886_ _0889_ _0847_ VGND VGND VPWR VPWR _0013_
+ sky130_fd_sc_hd__o211a_1
X_1398_ _0783_ _0789_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__or3b_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1321_ normal_mode_inst.timer_cnt\[7\] _0765_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nand2_1
X_1252_ phase_pwm_inst.counter\[22\] _0616_ _0718_ _0719_ VGND VGND VPWR VPWR _0194_
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1183_ phase_pwm_inst.counter\[16\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0660_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0967_ phase_pwm_inst.counter\[5\] VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__inv_2
X_1519_ _0925_ _0926_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1870_ net99 VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__inv_2
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1166_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__and2_1
X_1304_ _0635_ _0749_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__xnor2_1
X_1235_ _0707_ phase_pwm_inst.counter\[27\] _0616_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
X_1097_ phase_pwm_inst.counter\[13\] _0464_ _0567_ _0573_ _0569_ VGND VGND VPWR VPWR
+ _0574_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1020_ fast_pwm_inst.pwm_counter\[3\] VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__inv_2
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1922_ clknet_3_5__leaf_clk _0060_ _0105_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1784_ _0034_ _0420_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and2b_1
X_1853_ net99 VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__inv_2
X_1149_ _0624_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nand2_1
X_1218_ phase_pwm_inst.counter\[28\] _0470_ _0693_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or3b_1
XFILLER_20_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1003_ fast_pwm_inst.pwm_counter\[21\] VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__inv_2
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1905_ clknet_3_2__leaf_clk _0190_ _0088_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1767_ normal_mode_inst.timer_cnt\[19\] normal_mode_inst.timer_cnt\[20\] _0773_ normal_mode_inst.timer_cnt\[21\]
+ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__a31o_1
X_1836_ net99 VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__inv_2
XFILLER_1_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1698_ _0449_ net23 _0363_ _0364_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a221o_1
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1552_ _0477_ net50 _0919_ _0212_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a221o_1
X_1621_ _0446_ net60 net59 _0447_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__a22o_1
X_1483_ fast_pwm_inst.pwm_counter\[27\] _0898_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__and2_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1819_ net99 VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__inv_2
XFILLER_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0983_ net78 VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__inv_2
XFILLER_8_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1604_ fast_pwm_inst.pwm_counter\[27\] _0522_ _0523_ fast_pwm_inst.pwm_counter\[26\]
+ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o221a_1
X_1535_ _0941_ _0939_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__nand2b_1
X_1466_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__inv_2
X_1397_ net86 _0473_ _0474_ net85 _0782_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__o221a_1
XFILLER_37_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1320_ normal_mode_inst.timer_cnt\[5\] normal_mode_inst.timer_cnt\[4\] normal_mode_inst.timer_cnt\[6\]
+ _0763_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__and4_1
X_1182_ phase_pwm_inst.counter\[16\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0659_ sky130_fd_sc_hd__or2_1
X_1251_ _0677_ _0715_ _0616_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__o21ba_1
XFILLER_32_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0966_ phase_pwm_inst.counter\[6\] VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__inv_2
X_1518_ _0495_ net61 net60 _0496_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__a22o_1
X_1449_ _0876_ _0877_ _0847_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_2_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1303_ _0754_ phase_pwm_inst.counter\[6\] _0616_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1165_ phase_pwm_inst.counter\[8\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0642_
+ sky130_fd_sc_hd__xor2_1
X_1096_ _0566_ _0568_ _0552_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__a21boi_1
X_1234_ _0684_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__xor2_1
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0949_ phase_pwm_inst.counter\[24\] VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1852_ net99 VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__inv_2
X_1921_ clknet_3_5__leaf_clk _0049_ _0104_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1783_ normal_mode_inst.timer_cnt\[30\] _0780_ normal_mode_inst.timer_cnt\[31\] VGND
+ VGND VPWR VPWR _0420_ sky130_fd_sc_hd__a21o_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1079_ net76 phase_pwm_inst.counter\[1\] VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__and2b_1
X_1148_ phase_pwm_inst.counter\[1\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0625_
+ sky130_fd_sc_hd__or2_1
X_1217_ phase_pwm_inst.counter\[28\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0694_ sky130_fd_sc_hd__xor2_1
XFILLER_20_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1002_ fast_pwm_inst.pwm_counter\[22\] VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__inv_2
X_1835_ net99 VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__inv_2
X_1904_ clknet_3_2__leaf_clk _0189_ _0087_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_1766_ normal_mode_inst.timer_cnt\[20\] _0774_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__xnor2_1
X_1697_ phase_pwm_inst.counter\[3\] net26 VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__and2b_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1482_ fast_pwm_inst.pwm_counter\[27\] _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__or2_1
X_1551_ _0216_ _0217_ _0219_ _0221_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__or4_1
X_1620_ _0447_ net59 net58 _0448_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__o22a_1
XFILLER_39_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1818_ net99 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__inv_2
X_1749_ normal_mode_inst.timer_cnt\[10\] _0767_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_37_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0982_ net79 VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__inv_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1465_ fast_pwm_inst.pwm_counter\[21\] fast_pwm_inst.pwm_counter\[20\] fast_pwm_inst.pwm_counter\[19\]
+ _0882_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__and4_1
X_1603_ fast_pwm_inst.pwm_counter\[29\] _0520_ _0521_ fast_pwm_inst.pwm_counter\[28\]
+ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__o22a_1
X_1534_ _0936_ _0939_ _0941_ _0204_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or4_1
X_1396_ _0800_ _0835_ _0839_ _0804_ _0792_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__o32a_1
XFILLER_50_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1181_ phase_pwm_inst.direction _0614_ _0650_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a22o_1
X_1250_ _0677_ _0715_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nand2_1
XFILLER_32_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0965_ phase_pwm_inst.counter\[7\] VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__inv_2
X_1517_ _0496_ net60 net59 _0497_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__o22a_1
X_1448_ fast_pwm_inst.pwm_counter\[15\] _0874_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__or2_1
X_1379_ net66 _0491_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_24_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1302_ _0639_ _0751_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__xnor2_1
X_1233_ _0683_ _0687_ _0704_ _0682_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__o31a_1
X_1095_ phase_pwm_inst.counter\[8\] _0466_ _0570_ _0571_ VGND VGND VPWR VPWR _0572_
+ sky130_fd_sc_hd__o211a_1
X_1164_ phase_pwm_inst.direction _0604_ _0632_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__a22o_1
X_0948_ phase_pwm_inst.counter\[25\] VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1851_ net99 VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__inv_2
X_1920_ clknet_3_5__leaf_clk _0038_ _0103_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_1782_ normal_mode_inst.timer_cnt\[30\] _0780_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__xor2_1
XFILLER_6_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1216_ phase_pwm_inst.direction _0605_ _0680_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1078_ phase_pwm_inst.counter\[0\] net65 VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nand2b_1
X_1147_ phase_pwm_inst.counter\[1\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0624_
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1001_ fast_pwm_inst.pwm_counter\[23\] VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__inv_2
X_1765_ _0774_ _0413_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and2_1
X_1834_ net99 VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__inv_2
X_1903_ clknet_3_2__leaf_clk _0188_ _0086_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_1696_ _0449_ net23 net12 _0450_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_11_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1481_ _0898_ _0847_ _0897_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__and3b_1
X_1550_ fast_pwm_inst.pwm_counter\[24\] _0504_ _0220_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__o21ai_1
XFILLER_39_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1817_ net99 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__inv_2
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1748_ _0767_ _0406_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__and2b_1
X_1679_ _0342_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0981_ net80 VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__inv_2
X_1602_ _0268_ _0269_ _0270_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__or3b_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1464_ _0886_ _0887_ _0847_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__and3b_1
X_1395_ _0836_ _0837_ _0838_ _0801_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__or4b_1
X_1533_ fast_pwm_inst.pwm_counter\[11\] _0517_ _0935_ _0516_ fast_pwm_inst.pwm_counter\[12\]
+ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__o32ai_1
XFILLER_50_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1180_ _0656_ _0655_ _0654_ _0653_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__and4b_1
X_0964_ phase_pwm_inst.counter\[8\] VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__inv_2
X_1516_ _0497_ net59 _0920_ _0923_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__a221o_1
X_1378_ _0466_ fast_pwm_inst.pwm_counter\[8\] _0817_ _0821_ VGND VGND VPWR VPWR _0822_
+ sky130_fd_sc_hd__a31o_1
X_1447_ fast_pwm_inst.pwm_counter\[15\] fast_pwm_inst.pwm_counter\[14\] fast_pwm_inst.pwm_counter\[13\]
+ _0870_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and4_1
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1301_ _0753_ phase_pwm_inst.counter\[7\] _0616_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
X_1232_ _0687_ _0704_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__nor2_1
X_1094_ phase_pwm_inst.counter\[13\] _0464_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
X_1163_ _0635_ _0636_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__and3_1
X_0947_ phase_pwm_inst.counter\[26\] VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_30_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_41_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_44_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1781_ _0780_ _0419_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__nor2_1
X_1850_ net99 VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__inv_2
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1146_ phase_pwm_inst.counter\[2\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0623_
+ sky130_fd_sc_hd__and2_1
X_1215_ _0683_ _0684_ _0688_ _0691_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__or4bb_1
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1077_ phase_pwm_inst.counter\[1\] net76 VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nand2b_1
X_1979_ clknet_3_3__leaf_clk _0017_ _0162_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1000_ fast_pwm_inst.pwm_counter\[24\] VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__inv_2
X_1902_ clknet_3_0__leaf_clk _0187_ _0085_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[15\]
+ sky130_fd_sc_hd__dfrtp_2
X_1764_ normal_mode_inst.timer_cnt\[19\] _0773_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__or2_1
X_1833_ net99 VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__inv_2
X_1695_ _0450_ net12 net1 _0451_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a22o_1
X_1129_ _0601_ _0603_ _0604_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__or4_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1480_ fast_pwm_inst.pwm_counter\[26\] fast_pwm_inst.pwm_counter\[25\] _0893_ VGND
+ VGND VPWR VPWR _0898_ sky130_fd_sc_hd__and3_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1678_ phase_pwm_inst.counter\[27\] _0522_ _0523_ phase_pwm_inst.counter\[26\] _0345_
+ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__o221a_1
X_1816_ net99 VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__inv_2
X_1747_ normal_mode_inst.timer_cnt\[7\] normal_mode_inst.timer_cnt\[8\] _0765_ normal_mode_inst.timer_cnt\[9\]
+ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__a31o_1
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ net82 VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__inv_2
X_1601_ fast_pwm_inst.pwm_counter\[25\] _0524_ _0525_ fast_pwm_inst.pwm_counter\[24\]
+ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__a22o_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1532_ fast_pwm_inst.pwm_counter\[14\] _0514_ _0937_ _0940_ VGND VGND VPWR VPWR _0941_
+ sky130_fd_sc_hd__a211o_1
X_1463_ _0482_ _0884_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__nand2_1
X_1394_ _0461_ fast_pwm_inst.pwm_counter\[21\] _0792_ _0793_ VGND VGND VPWR VPWR _0838_
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0963_ phase_pwm_inst.counter\[9\] VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__inv_2
X_1515_ fast_pwm_inst.pwm_counter\[3\] _0519_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nor2_1
X_1377_ net67 _0490_ _0491_ net66 VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__a22o_1
X_1446_ _0874_ _0875_ _0847_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__and3b_1
XFILLER_23_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_48_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1162_ _0637_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__nor2_1
X_1300_ _0636_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__xnor2_1
X_1231_ _0680_ _0689_ _0690_ _0685_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__o211a_1
X_1093_ _0444_ net94 _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__a21oi_1
X_0946_ phase_pwm_inst.counter\[27\] VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__inv_2
XFILLER_9_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1429_ fast_pwm_inst.pwm_counter\[9\] fast_pwm_inst.pwm_counter\[8\] fast_pwm_inst.pwm_counter\[7\]
+ _0858_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__and4_1
XFILLER_28_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ normal_mode_inst.timer_cnt\[28\] _0779_ normal_mode_inst.timer_cnt\[29\] VGND
+ VGND VPWR VPWR _0419_ sky130_fd_sc_hd__a21oi_1
XFILLER_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1145_ _0448_ _0470_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__nor2_1
X_1214_ _0689_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_50_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1076_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__inv_2
X_1978_ clknet_3_3__leaf_clk _0016_ _0161_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_20_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1832_ net99 VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__inv_2
X_1901_ clknet_3_0__leaf_clk _0186_ _0084_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[14\]
+ sky130_fd_sc_hd__dfrtp_4
X_1763_ _0773_ _0412_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and2b_1
X_1694_ net26 phase_pwm_inst.counter\[3\] VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__nand2b_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1059_ net99 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
XFILLER_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1128_ phase_pwm_inst.counter\[27\] phase_pwm_inst.counter\[26\] phase_pwm_inst.counter\[25\]
+ phase_pwm_inst.counter\[24\] VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or4_1
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1815_ net99 VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__inv_2
XFILLER_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1677_ phase_pwm_inst.counter\[24\] _0525_ _0344_ _0343_ VGND VGND VPWR VPWR _0345_
+ sky130_fd_sc_hd__a31o_1
X_1746_ normal_mode_inst.timer_cnt\[8\] _0766_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__xnor2_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1462_ _0482_ _0884_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nor2_1
X_1600_ _0472_ net24 net22 _0473_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__o22a_1
X_1531_ _0487_ net38 net37 _0488_ _0938_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__a221o_1
X_1393_ _0794_ _0796_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nand2_1
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1729_ _0425_ net20 net19 _0426_ _0342_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0962_ phase_pwm_inst.counter\[10\] VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__inv_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ _0499_ net55 _0921_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__a22o_1
X_1445_ _0487_ _0872_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__nand2_1
X_1376_ net96 _0492_ _0816_ _0818_ _0819_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__o221a_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1230_ _0680_ _0689_ _0690_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__o21a_1
X_1092_ _0439_ net68 VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_1
X_1161_ phase_pwm_inst.counter\[6\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0638_
+ sky130_fd_sc_hd__nor2_1
X_0945_ phase_pwm_inst.counter\[28\] VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__inv_2
XFILLER_9_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1428_ _0862_ _0863_ _0847_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and3b_1
X_1359_ _0795_ _0802_ _0461_ fast_pwm_inst.pwm_counter\[21\] VGND VGND VPWR VPWR _0803_
+ sky130_fd_sc_hd__a2bb2o_1
Xclkload2 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_8
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ phase_pwm_inst.counter\[24\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0690_ sky130_fd_sc_hd__nand2_1
XFILLER_37_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1075_ _0439_ net68 _0465_ phase_pwm_inst.counter\[11\] VGND VGND VPWR VPWR _0552_
+ sky130_fd_sc_hd__o2bb2a_1
X_1144_ phase_pwm_inst.counter\[3\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0621_
+ sky130_fd_sc_hd__or2_1
X_1977_ clknet_3_3__leaf_clk _0015_ _0160_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1831_ net99 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__inv_2
X_1900_ clknet_3_0__leaf_clk _0185_ _0083_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_1762_ normal_mode_inst.timer_cnt\[17\] normal_mode_inst.timer_cnt\[16\] _0771_ normal_mode_inst.timer_cnt\[18\]
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a31o_1
X_1693_ _0430_ net15 _0351_ _0358_ _0359_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o221a_1
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1058_ net2 VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__inv_2
X_1127_ phase_pwm_inst.counter\[7\] phase_pwm_inst.counter\[6\] phase_pwm_inst.counter\[5\]
+ phase_pwm_inst.counter\[4\] VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__or4_1
XFILLER_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1814_ net99 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1745_ _0766_ _0405_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__and2_1
X_1676_ _0427_ net18 VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nand2_1
XFILLER_7_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1461_ _0847_ _0884_ _0885_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__and3_1
X_1392_ net72 _0486_ _0795_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a21o_1
X_1530_ fast_pwm_inst.pwm_counter\[13\] _0515_ _0516_ fast_pwm_inst.pwm_counter\[12\]
+ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__a22o_1
X_1728_ _0427_ net18 net17 _0428_ _0340_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__a221o_1
X_1659_ _0425_ net52 net51 _0426_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_5_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0961_ phase_pwm_inst.counter\[11\] VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1513_ _0499_ net55 net44 _0500_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__o22a_1
X_1375_ _0466_ fast_pwm_inst.pwm_counter\[8\] VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__nand2_1
X_1444_ _0487_ _0872_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1091_ _0441_ net66 net96 _0442_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a22o_1
X_1160_ _0445_ _0470_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__nor2_1
X_0944_ phase_pwm_inst.counter\[29\] VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__inv_2
X_1358_ _0797_ _0798_ _0800_ _0796_ _0801_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_38_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1427_ _0493_ _0860_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nand2_1
XFILLER_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1289_ _0745_ phase_pwm_inst.counter\[11\] _0616_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XFILLER_50_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload3 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__inv_12
XPHY_EDGE_ROW_3_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1212_ phase_pwm_inst.counter\[24\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0689_ sky130_fd_sc_hd__nor2_1
X_1143_ phase_pwm_inst.counter\[3\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0620_
+ sky130_fd_sc_hd__nor2_1
X_1074_ _0438_ net70 VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__nand2_1
X_1976_ clknet_3_3__leaf_clk _0014_ _0159_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_45_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1761_ normal_mode_inst.timer_cnt\[17\] _0772_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__xnor2_1
X_1830_ net99 VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__inv_2
X_1692_ _0430_ net15 VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__nor2_1
X_1126_ phase_pwm_inst.counter\[31\] phase_pwm_inst.counter\[28\] _0602_ VGND VGND
+ VPWR VPWR _0603_ sky130_fd_sc_hd__or3_1
X_1057_ net4 VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__inv_2
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1959_ clknet_3_4__leaf_clk _0027_ _0142_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1744_ normal_mode_inst.timer_cnt\[7\] _0765_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__or2_1
X_1813_ net99 VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__inv_2
X_1675_ phase_pwm_inst.counter\[26\] _0523_ _0524_ phase_pwm_inst.counter\[25\] VGND
+ VGND VPWR VPWR _0343_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1109_ phase_pwm_inst.counter\[25\] _0458_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1460_ fast_pwm_inst.pwm_counter\[19\] _0882_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__or2_1
X_1391_ _0829_ _0831_ _0833_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__o211a_1
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1658_ _0323_ _0324_ _0325_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__or4_1
X_1727_ _0350_ _0361_ _0391_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__o22a_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1589_ _0252_ _0256_ _0257_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_5_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0960_ phase_pwm_inst.counter\[12\] VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__inv_2
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1512_ _0500_ net44 net33 _0501_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1374_ net95 _0493_ _0494_ net94 _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a221o_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1443_ _0847_ _0872_ _0873_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1090_ _0442_ net96 net95 _0443_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__o221ai_2
X_0943_ phase_pwm_inst.counter\[30\] VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__inv_2
X_1357_ net77 _0482_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1426_ _0493_ _0860_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__nor2_1
X_1288_ _0648_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__xnor2_1
XFILLER_18_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload4 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_8
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1142_ _0617_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__nor2_1
X_1211_ _0686_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__nor2_1
X_1073_ _0539_ _0549_ _0538_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__a21o_1
X_1975_ clknet_3_2__leaf_clk _0013_ _0158_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_29_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1409_ _0499_ _0848_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nor2_1
XFILLER_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1760_ _0772_ _0411_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__and2_1
X_1691_ _0429_ net16 net14 _0431_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__o22a_1
X_1125_ phase_pwm_inst.counter\[30\] phase_pwm_inst.counter\[29\] VGND VGND VPWR VPWR
+ _0602_ sky130_fd_sc_hd__or2_1
X_1056_ net5 VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__inv_2
X_1958_ clknet_3_4__leaf_clk _0026_ _0141_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1889_ clknet_3_4__leaf_clk _0174_ _0072_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1674_ phase_pwm_inst.counter\[28\] _0521_ _0522_ phase_pwm_inst.counter\[27\] VGND
+ VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a22o_1
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1812_ net99 VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__inv_2
X_1743_ _0765_ _0404_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__and2b_1
X_1108_ _0423_ net86 net85 _0424_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__a22o_1
X_1039_ net35 VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__inv_2
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1390_ net70 _0487_ _0827_ _0825_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__o31a_1
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1588_ fast_pwm_inst.pwm_counter\[20\] _0527_ _0528_ fast_pwm_inst.pwm_counter\[19\]
+ _0253_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__a221o_1
X_1726_ _0353_ _0356_ _0392_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or4_1
X_1657_ _0422_ net56 net54 _0423_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o22ai_1
XFILLER_7_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1511_ fast_pwm_inst.pwm_counter\[3\] _0519_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1442_ fast_pwm_inst.pwm_counter\[13\] _0870_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2_1
X_1373_ net96 _0492_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__and2_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1709_ phase_pwm_inst.counter\[10\] _0536_ _0375_ _0376_ VGND VGND VPWR VPWR _0377_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_24_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0942_ phase_pwm_inst.counter\[31\] VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__inv_2
X_1425_ _0847_ _0860_ _0861_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__and3_1
X_1356_ _0798_ _0799_ _0797_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_38_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1287_ phase_pwm_inst.counter\[10\] phase_pwm_inst.direction _0743_ VGND VGND VPWR
+ VPWR _0744_ sky130_fd_sc_hd__a21oi_1
Xclkload5 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_4
XFILLER_10_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1072_ _0542_ _0544_ _0545_ _0546_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a311o_1
X_1141_ phase_pwm_inst.counter\[4\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0618_
+ sky130_fd_sc_hd__nor2_1
X_1210_ phase_pwm_inst.counter\[25\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0687_ sky130_fd_sc_hd__nor2_1
XFILLER_45_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1974_ clknet_3_2__leaf_clk _0012_ _0157_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1408_ _0499_ _0848_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__nand2_1
XFILLER_45_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1339_ _0457_ fast_pwm_inst.pwm_counter\[26\] fast_pwm_inst.pwm_counter\[25\] _0458_
+ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a22o_1
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1690_ _0432_ net13 _0354_ _0355_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o221a_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1124_ phase_pwm_inst.counter\[3\] phase_pwm_inst.counter\[2\] phase_pwm_inst.counter\[1\]
+ phase_pwm_inst.counter\[0\] VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__or4_1
X_1055_ net6 VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__inv_2
X_1957_ clknet_3_4__leaf_clk _0025_ _0140_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_1888_ clknet_3_4__leaf_clk _0173_ _0071_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1811_ net99 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__inv_2
X_1673_ phase_pwm_inst.counter\[29\] _0520_ _0521_ phase_pwm_inst.counter\[28\] VGND
+ VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o22a_1
XFILLER_7_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1742_ normal_mode_inst.timer_cnt\[5\] normal_mode_inst.timer_cnt\[4\] _0763_ normal_mode_inst.timer_cnt\[6\]
+ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__a31o_1
X_1107_ _0537_ _0550_ _0579_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1038_ net36 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__inv_2
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1725_ phase_pwm_inst.counter\[20\] _0527_ net8 _0436_ _0360_ VGND VGND VPWR VPWR
+ _0393_ sky130_fd_sc_hd__a221o_1
X_1587_ fast_pwm_inst.pwm_counter\[21\] _0526_ net8 _0486_ _0254_ VGND VGND VPWR VPWR
+ _0257_ sky130_fd_sc_hd__a221o_1
X_1656_ _0421_ net57 net56 _0422_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__a22o_1
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1510_ _0909_ _0918_ _0479_ net48 VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1441_ fast_pwm_inst.pwm_counter\[13\] _0870_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__nand2_1
X_1372_ net94 _0494_ _0813_ _0814_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_33_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1708_ _0440_ net3 VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and2_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1639_ phase_pwm_inst.counter\[23\] _0505_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nor2_1
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_50_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1355_ net74 _0484_ _0485_ net73 VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a22o_1
X_1424_ fast_pwm_inst.pwm_counter\[7\] _0858_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_38_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1286_ _0742_ _0644_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2b_1
XFILLER_50_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload6 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1071_ _0543_ _0547_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__nor2_1
X_1140_ _0447_ _0470_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__nor2_1
X_1973_ clknet_3_2__leaf_clk _0010_ _0156_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_2
X_1338_ _0456_ fast_pwm_inst.pwm_counter\[27\] fast_pwm_inst.pwm_counter\[26\] _0457_
+ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__o22a_1
X_1407_ _0847_ _0848_ _0849_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__and3_1
XFILLER_51_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1269_ phase_pwm_inst.counter\[16\] _0616_ _0662_ _0730_ VGND VGND VPWR VPWR _0188_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_7_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1123_ _0595_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__or2_1
X_1054_ net7 VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__inv_2
X_1956_ clknet_3_4__leaf_clk _0022_ _0139_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_1887_ clknet_3_4__leaf_clk _0172_ _0070_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ net99 VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__inv_2
XFILLER_15_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1741_ normal_mode_inst.timer_cnt\[5\] _0764_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__xnor2_1
X_1672_ _0422_ net24 _0520_ phase_pwm_inst.counter\[29\] VGND VGND VPWR VPWR _0340_
+ sky130_fd_sc_hd__a2bb2o_1
X_1106_ _0541_ _0544_ _0547_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__and4b_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1037_ net37 VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__inv_2
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1939_ clknet_3_7__leaf_clk _0048_ _0122_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput90 TIMER_TOP[3] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_44_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1724_ _0349_ _0351_ _0352_ _0359_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__or4b_1
X_1586_ fast_pwm_inst.pwm_counter\[17\] _0530_ _0531_ fast_pwm_inst.pwm_counter\[16\]
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__a22o_1
X_1655_ phase_pwm_inst.counter\[25\] _0503_ _0504_ phase_pwm_inst.counter\[24\] VGND
+ VGND VPWR VPWR _0324_ sky130_fd_sc_hd__a22o_1
XFILLER_41_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_36_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1371_ _0467_ fast_pwm_inst.pwm_counter\[6\] VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nand2_1
XFILLER_4_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1440_ _0870_ _0871_ _0847_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_33_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1638_ _0434_ net42 net41 _0435_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a221o_1
X_1707_ _0441_ net2 net32 _0442_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__a22o_1
X_1569_ _0495_ net29 net28 _0496_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_1
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1354_ net75 _0483_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and2_1
X_1423_ fast_pwm_inst.pwm_counter\[7\] _0858_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__nand2_1
X_1285_ _0645_ _0741_ _0646_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__o21ai_1
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1070_ _0432_ net77 net75 _0433_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o22a_1
X_1972_ clknet_3_2__leaf_clk _0009_ _0155_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_23_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1337_ _0453_ fast_pwm_inst.pwm_counter\[30\] fast_pwm_inst.pwm_counter\[29\] _0454_
+ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__o22a_1
X_1406_ fast_pwm_inst.pwm_counter\[1\] fast_pwm_inst.pwm_counter\[0\] VGND VGND VPWR
+ VPWR _0849_ sky130_fd_sc_hd__or2_1
X_1268_ _0616_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__nor2_1
XFILLER_51_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1199_ _0674_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__nand2b_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1122_ _0421_ net89 _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__o21ai_1
X_1053_ net8 VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__inv_2
XFILLER_18_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1955_ clknet_3_5__leaf_clk _0011_ _0138_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_1886_ net99 VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__inv_2
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0421_ net25 net24 _0422_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__a22o_1
X_1740_ _0764_ _0403_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__and2_1
X_1105_ _0538_ _0539_ _0580_ _0581_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_16_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1036_ net38 VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__inv_2
X_1869_ net99 VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
X_1938_ clknet_3_7__leaf_clk _0047_ _0121_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[18\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput91 TIMER_TOP[4] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput80 TIMER_TOP[23] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1654_ _0423_ net54 net53 _0424_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__a22o_1
X_1723_ _0381_ _0388_ _0389_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__and4b_1
X_1585_ _0485_ net9 VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__nand2_1
XFILLER_41_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1019_ fast_pwm_inst.pwm_counter\[4\] VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1370_ net93 _0495_ _0496_ net92 VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__a22o_1
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1637_ _0432_ net45 net43 _0433_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__a221o_1
X_1706_ _0371_ _0372_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o21a_1
XFILLER_48_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1499_ phase_pwm_inst.pwm_outa _0907_ _0908_ fast_pwm_inst.pwm_outa VGND VGND VPWR
+ VPWR net100 sky130_fd_sc_hd__a22o_2
X_1568_ _0497_ net27 net26 _0498_ _0237_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__a221o_1
XFILLER_14_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ _0858_ _0859_ _0847_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__and3b_1
X_1353_ net75 _0483_ _0484_ net74 VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__o22a_1
X_1284_ phase_pwm_inst.counter\[8\] phase_pwm_inst.direction _0643_ VGND VGND VPWR
+ VPWR _0741_ sky130_fd_sc_hd__a21o_1
X_0999_ fast_pwm_inst.pwm_counter\[25\] VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1971_ clknet_3_2__leaf_clk _0008_ _0154_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_1405_ fast_pwm_inst.pwm_counter\[1\] fast_pwm_inst.pwm_counter\[0\] VGND VGND VPWR
+ VPWR _0848_ sky130_fd_sc_hd__nand2_1
Xinput1 PWM_CNTA[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_1336_ normal_mode_inst.timer_cnt\[30\] normal_mode_inst.timer_cnt\[31\] _0780_ VGND
+ VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and3_1
XFILLER_36_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1198_ phase_pwm_inst.counter\[21\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0675_ sky130_fd_sc_hd__or2_1
X_1267_ _0658_ _0661_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__and2b_1
XFILLER_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1052_ net9 VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__inv_2
X_1121_ _0585_ _0593_ _0594_ _0597_ _0588_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__a221o_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1954_ clknet_3_5__leaf_clk _0000_ _0137_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1885_ net99 VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__inv_2
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1319_ normal_mode_inst.timer_cnt\[4\] _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__nand2_1
XFILLER_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1670_ _0421_ net57 _0325_ _0338_ _0334_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__o221a_1
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1104_ _0436_ net72 _0537_ _0540_ _0545_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__o2111a_1
X_1035_ net39 VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__inv_2
X_1937_ clknet_3_6__leaf_clk _0046_ _0120_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput81 TIMER_TOP[24] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
Xinput70 TIMER_TOP[14] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_2
X_1868_ net99 VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__inv_2
Xinput92 TIMER_TOP[5] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlymetal6s2s_1
X_1799_ net99 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__inv_2
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ fast_pwm_inst.pwm_counter\[20\] _0527_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__nor2_1
X_1653_ _0304_ _0315_ _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a21oi_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1722_ net6 _0383_ phase_pwm_inst.counter\[14\] VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or3b_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1018_ fast_pwm_inst.pwm_counter\[5\] VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1705_ _0442_ net32 net31 _0443_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__o22a_1
X_1636_ phase_pwm_inst.counter\[21\] _0507_ _0508_ phase_pwm_inst.counter\[20\] VGND
+ VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a22o_1
X_1567_ _0498_ net26 _0234_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__o22a_1
X_1498_ phase_pwm_inst.pwm_outb _0907_ _0908_ fast_pwm_inst.pwm_outb VGND VGND VPWR
+ VPWR net101 sky130_fd_sc_hd__a22o_1
XFILLER_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1421_ fast_pwm_inst.pwm_counter\[6\] _0856_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or2_1
XFILLER_48_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1352_ net73 _0485_ _0486_ net72 VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__o22a_1
X_1283_ _0740_ phase_pwm_inst.counter\[12\] _0616_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ fast_pwm_inst.pwm_counter\[26\] VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__inv_2
X_1619_ _0285_ _0286_ _0287_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21o_1
XFILLER_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1970_ clknet_3_2__leaf_clk _0007_ _0153_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_1335_ normal_mode_inst.timer_cnt\[29\] normal_mode_inst.timer_cnt\[28\] _0779_ VGND
+ VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and3_1
XFILLER_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1404_ _0501_ _0847_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__and2_1
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 PWM_CNTA[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
X_1266_ _0728_ phase_pwm_inst.counter\[17\] _0616_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
X_1197_ _0431_ _0470_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__nor2_1
XFILLER_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1051_ net10 VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__inv_2
X_1120_ _0589_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__nand2_1
X_1953_ clknet_3_6__leaf_clk _0032_ _0136_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_outa
+ sky130_fd_sc_hd__dfrtp_1
X_1884_ net99 VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__inv_2
X_1318_ normal_mode_inst.timer_cnt\[0\] normal_mode_inst.timer_cnt\[1\] normal_mode_inst.timer_cnt\[3\]
+ normal_mode_inst.timer_cnt\[2\] VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__and4_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1249_ _0717_ phase_pwm_inst.counter\[23\] _0616_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1034_ net40 VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__inv_2
X_1103_ _0436_ net72 net71 _0437_ _0546_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__a221oi_1
X_1936_ clknet_3_7__leaf_clk _0045_ _0119_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_1867_ net99 VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__inv_2
Xinput60 PWM_CNTB[5] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
Xinput71 TIMER_TOP[15] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput82 TIMER_TOP[25] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
Xinput93 TIMER_TOP[6] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
X_1798_ net99 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1721_ _0386_ _0384_ _0385_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or3b_1
X_1583_ _0483_ net11 net10 _0484_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__a22o_1
X_1652_ _0309_ _0320_ _0316_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_36_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ fast_pwm_inst.pwm_counter\[6\] VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__inv_2
X_1919_ clknet_3_6__leaf_clk _0034_ _0102_ VGND VGND VPWR VPWR irq_timer_normal sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1704_ _0443_ net31 net30 _0444_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a22o_1
X_1497_ net98 net97 VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__and2b_1
X_1566_ _0499_ net23 net12 _0500_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o221a_1
X_1635_ _0437_ net39 net38 _0438_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__o221ai_2
XTAP_TAPCELL_ROW_32_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1351_ net77 _0482_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__and2_1
X_1420_ fast_pwm_inst.pwm_counter\[6\] fast_pwm_inst.pwm_counter\[5\] fast_pwm_inst.pwm_counter\[4\]
+ _0852_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__and4_1
XFILLER_48_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1282_ _0731_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_21_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0997_ fast_pwm_inst.pwm_counter\[27\] VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__inv_2
X_1618_ _0448_ net58 net55 _0449_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a22o_1
X_1549_ _0476_ net51 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2_1
XFILLER_5_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1334_ normal_mode_inst.timer_cnt\[27\] _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__and2_1
X_1403_ _0790_ _0791_ _0840_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o22a_4
X_1265_ _0666_ _0722_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__xnor2_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 PWM_CNTA[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
X_1196_ _0671_ _0672_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__nand2_1
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1050_ net11 VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__inv_2
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1883_ net99 VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
X_1952_ clknet_3_6__leaf_clk _0033_ _0135_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_outb
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1317_ normal_mode_inst.timer_cnt\[0\] normal_mode_inst.timer_cnt\[1\] normal_mode_inst.timer_cnt\[2\]
+ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__and3_1
X_1248_ _0672_ _0716_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__xor2_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1179_ phase_pwm_inst.counter\[15\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0656_ sky130_fd_sc_hd__xnor2_1
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1102_ _0551_ _0577_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__a21bo_1
X_1033_ net41 VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__inv_2
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 PWM_CNTB[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput72 TIMER_TOP[16] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
X_1935_ clknet_3_7__leaf_clk _0044_ _0118_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[15\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput61 PWM_CNTB[6] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
X_1797_ net99 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__inv_2
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1866_ net99 VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__inv_2
Xinput94 TIMER_TOP[7] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
Xinput83 TIMER_TOP[26] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1651_ _0305_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__nor2_1
X_1720_ _0380_ _0384_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_13_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1582_ _0480_ net15 net14 _0481_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a22o_1
X_1016_ fast_pwm_inst.pwm_counter\[7\] VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_14_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1849_ net99 VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__inv_2
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1918_ clknet_3_5__leaf_clk _0203_ _0101_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1703_ _0444_ net30 net29 _0445_ _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o221a_1
X_1634_ _0438_ net38 _0283_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__a22o_1
X_1496_ net97 net98 VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and2b_1
X_1565_ _0500_ net12 net1 _0501_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1350_ _0460_ fast_pwm_inst.pwm_counter\[22\] fast_pwm_inst.pwm_counter\[21\] _0461_
+ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__o22a_1
X_1281_ _0612_ _0650_ _0655_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__nor3_1
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0996_ fast_pwm_inst.pwm_counter\[28\] VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__inv_2
XFILLER_5_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1617_ _0449_ net55 net44 _0450_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__o22a_1
X_1479_ fast_pwm_inst.pwm_counter\[26\] _0896_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or2_1
X_1548_ _0473_ net54 net53 _0474_ _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a221o_1
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1402_ _0842_ _0844_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__or3b_1
XFILLER_5_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 PWM_CNTA[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
X_1333_ normal_mode_inst.timer_cnt\[25\] normal_mode_inst.timer_cnt\[26\] _0777_ VGND
+ VGND VPWR VPWR _0778_ sky130_fd_sc_hd__and3_1
X_1264_ _0724_ _0727_ phase_pwm_inst.counter\[18\] _0616_ VGND VGND VPWR VPWR _0190_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1195_ phase_pwm_inst.counter\[23\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0672_ sky130_fd_sc_hd__xor2_1
X_0979_ net83 VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__inv_2
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1882_ net99 VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__inv_2
X_1951_ clknet_3_6__leaf_clk _0062_ _0134_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1178_ phase_pwm_inst.counter\[12\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0655_ sky130_fd_sc_hd__xor2_1
X_1316_ phase_pwm_inst.counter\[0\] _0616_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__xnor2_1
X_1247_ _0675_ _0678_ _0714_ phase_pwm_inst.direction phase_pwm_inst.counter\[22\]
+ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_44_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1032_ net42 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__inv_2
X_1101_ _0437_ net71 net70 _0438_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__o22a_1
XFILLER_46_271 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1934_ clknet_3_7__leaf_clk _0043_ _0117_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput84 TIMER_TOP[27] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
Xinput40 PWM_CNTB[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_1
X_1796_ net99 VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_2
Xinput51 PWM_CNTB[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput62 PWM_CNTB[7] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 TIMER_TOP[17] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput95 TIMER_TOP[8] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
X_1865_ net99 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__inv_2
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1650_ phase_pwm_inst.counter\[20\] _0508_ _0509_ phase_pwm_inst.counter\[19\] _0318_
+ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o221a_1
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1581_ _0228_ _0233_ _0248_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o22a_1
XFILLER_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1015_ fast_pwm_inst.pwm_counter\[8\] VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__inv_2
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1917_ clknet_3_7__leaf_clk _0202_ _0100_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_1779_ normal_mode_inst.timer_cnt\[28\] _0779_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__xor2_1
X_1848_ net99 VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1564_ _0499_ net23 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__and2_1
X_1702_ _0367_ _0368_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21o_1
X_1633_ _0298_ _0299_ _0301_ _0282_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_1_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _0470_ _0600_ _0615_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__a21o_1
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1280_ _0738_ phase_pwm_inst.counter\[13\] _0616_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux2_1
XFILLER_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0995_ fast_pwm_inst.pwm_counter\[29\] VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__inv_2
X_1547_ _0471_ net57 net56 _0472_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a22o_1
X_1616_ _0450_ net44 net33 _0451_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a22o_1
X_1478_ _0896_ _0847_ _0895_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__and3b_1
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1401_ _0458_ fast_pwm_inst.pwm_counter\[25\] _0478_ net81 _0781_ VGND VGND VPWR
+ VPWR _0845_ sky130_fd_sc_hd__o221a_1
XFILLER_5_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 PWM_CNTA[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
X_1332_ normal_mode_inst.timer_cnt\[23\] normal_mode_inst.timer_cnt\[22\] normal_mode_inst.timer_cnt\[24\]
+ _0775_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__and4_1
X_1263_ _0663_ _0668_ _0723_ _0616_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__a31o_1
X_1194_ phase_pwm_inst.counter\[20\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0671_ sky130_fd_sc_hd__xor2_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0978_ net84 VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__inv_2
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1950_ clknet_3_7__leaf_clk _0061_ _0133_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1881_ net99 VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__inv_2
X_1315_ _0761_ phase_pwm_inst.counter\[1\] _0616_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1177_ phase_pwm_inst.counter\[14\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0654_ sky130_fd_sc_hd__xor2_1
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1246_ _0675_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__nand2_1
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1031_ net43 VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__inv_2
X_1100_ _0565_ _0572_ _0576_ _0575_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__a31o_1
X_1933_ clknet_3_7__leaf_clk _0042_ _0116_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput96 TIMER_TOP[9] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_2
Xinput85 TIMER_TOP[28] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
Xinput52 PWM_CNTB[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
Xinput74 TIMER_TOP[18] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 PWM_CNTB[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
X_1795_ net99 VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__inv_2
Xinput30 PWM_CNTA[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput63 PWM_CNTB[8] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_1
X_1864_ net99 VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__inv_2
X_1229_ _0702_ phase_pwm_inst.counter\[28\] _0616_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1580_ _0229_ _0231_ _0232_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__or4_1
XFILLER_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1014_ fast_pwm_inst.pwm_counter\[9\] VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__inv_2
XFILLER_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1847_ net99 VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__inv_2
X_1916_ clknet_3_7__leaf_clk _0201_ _0099_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_1778_ _0779_ _0418_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__nor2_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1701_ _0445_ net29 net28 _0446_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__a22o_1
X_1494_ _0471_ _0906_ _0847_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__a21boi_1
X_1632_ phase_pwm_inst.counter\[11\] _0517_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__o21ai_1
X_1563_ _0230_ _0232_ _0229_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_1_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0994_ fast_pwm_inst.pwm_counter\[30\] VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__inv_2
X_1477_ _0477_ _0894_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nor2_1
X_1546_ _0213_ _0214_ _0215_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__or3b_1
X_1615_ _0446_ net60 VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or2_1
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1400_ net81 _0478_ _0791_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__a211o_1
X_1331_ normal_mode_inst.timer_cnt\[22\] _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nand2_1
XFILLER_5_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1262_ _0726_ phase_pwm_inst.counter\[19\] _0616_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
Xinput6 PWM_CNTA[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
X_1193_ _0661_ _0669_ _0658_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__nand3b_1
X_0977_ net85 VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__inv_2
X_1529_ fast_pwm_inst.pwm_counter\[15\] _0513_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nor2_1
XFILLER_42_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1880_ net99 VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1314_ phase_pwm_inst.counter\[0\] _0626_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1176_ _0651_ _0652_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__and2b_1
X_1245_ phase_pwm_inst.counter\[20\] phase_pwm_inst.direction _0674_ _0712_ VGND VGND
+ VPWR VPWR _0714_ sky130_fd_sc_hd__a211o_1
XFILLER_7_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1030_ net45 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__inv_2
X_1932_ clknet_3_7__leaf_clk _0041_ _0115_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput20 PWM_CNTA[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 PWM_CNTA[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1863_ net99 VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
Xinput97 TMR_MODE[0] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
X_1794_ net99 VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_2
Xinput42 PWM_CNTB[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
Xinput64 PWM_CNTB[9] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput53 PWM_CNTB[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput86 TIMER_TOP[29] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
Xinput75 TIMER_TOP[19] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1228_ _0693_ _0694_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1159_ phase_pwm_inst.counter\[7\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0636_
+ sky130_fd_sc_hd__xor2_1
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1013_ fast_pwm_inst.pwm_counter\[10\] VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__inv_2
X_1777_ normal_mode_inst.timer_cnt\[27\] _0778_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor2_1
X_1846_ net99 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__inv_2
X_1915_ clknet_3_5__leaf_clk _0200_ _0098_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1700_ _0446_ net28 net27 _0447_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o22a_1
X_1631_ phase_pwm_inst.counter\[13\] _0515_ _0516_ phase_pwm_inst.counter\[12\] VGND
+ VGND VPWR VPWR _0300_ sky130_fd_sc_hd__o22a_1
X_1493_ _0847_ _0905_ _0906_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__and3_1
X_1562_ fast_pwm_inst.pwm_counter\[13\] _0534_ _0535_ fast_pwm_inst.pwm_counter\[12\]
+ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1829_ net99 VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__inv_2
XFILLER_38_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0993_ fast_pwm_inst.pwm_counter\[31\] VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__inv_2
X_1614_ phase_pwm_inst.counter\[13\] _0515_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__o21ai_1
X_1476_ fast_pwm_inst.pwm_counter\[25\] _0893_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__or2_1
XFILLER_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1545_ fast_pwm_inst.pwm_counter\[25\] _0503_ _0504_ fast_pwm_inst.pwm_counter\[24\]
+ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1330_ normal_mode_inst.timer_cnt\[19\] normal_mode_inst.timer_cnt\[21\] normal_mode_inst.timer_cnt\[20\]
+ _0773_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__and4_1
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1261_ _0667_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__xnor2_1
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1192_ _0668_ _0667_ _0665_ _0663_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__and4b_1
Xinput7 PWM_CNTA[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0976_ net86 VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__inv_2
XFILLER_10_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1459_ fast_pwm_inst.pwm_counter\[19\] _0882_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__nand2_1
X_1528_ fast_pwm_inst.pwm_counter\[15\] _0513_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__and2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1313_ _0760_ phase_pwm_inst.counter\[2\] _0616_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
X_1244_ phase_pwm_inst.counter\[20\] phase_pwm_inst.direction _0712_ VGND VGND VPWR
+ VPWR _0713_ sky130_fd_sc_hd__a21o_1
X_1175_ phase_pwm_inst.counter\[13\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0652_ sky130_fd_sc_hd__or2_1
X_0959_ phase_pwm_inst.counter\[14\] VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__inv_2
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1931_ clknet_3_7__leaf_clk _0040_ _0114_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput32 PWM_CNTA[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 PWM_CNTB[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__buf_1
Xinput21 PWM_CNTA[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput54 PWM_CNTB[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_1793_ net99 VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__inv_2
X_1862_ net99 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__inv_2
Xinput10 PWM_CNTA[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
Xinput87 TIMER_TOP[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
Xinput98 TMR_MODE[1] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
Xinput76 TIMER_TOP[1] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
Xinput65 TIMER_TOP[0] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_1
X_1227_ _0423_ _0701_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__xnor2_1
X_1158_ _0633_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__nor2_1
X_1089_ _0440_ net67 net66 _0441_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__o22a_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_7_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1012_ fast_pwm_inst.pwm_counter\[11\] VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__inv_2
XFILLER_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1914_ clknet_3_4__leaf_clk _0199_ _0097_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_1845_ net99 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__inv_2
X_1776_ _0778_ _0417_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__nor2_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1630_ _0440_ net35 net34 _0441_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o22a_1
X_1492_ fast_pwm_inst.pwm_counter\[30\] _0904_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nand2_1
X_1561_ _0487_ net6 net5 _0488_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1759_ normal_mode_inst.timer_cnt\[16\] _0771_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or2_1
X_1828_ net99 VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__inv_2
XFILLER_13_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0992_ phase_pwm_inst.direction VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__inv_2
X_1544_ _0472_ net56 net54 _0473_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o22a_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1613_ phase_pwm_inst.counter\[13\] _0515_ _0516_ phase_pwm_inst.counter\[12\] VGND
+ VGND VPWR VPWR _0282_ sky130_fd_sc_hd__a22o_1
X_1475_ fast_pwm_inst.pwm_counter\[24\] _0891_ _0894_ _0847_ VGND VGND VPWR VPWR _0016_
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 PWM_CNTA[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
X_1260_ phase_pwm_inst.counter\[18\] phase_pwm_inst.direction _0724_ VGND VGND VPWR
+ VPWR _0725_ sky130_fd_sc_hd__a21oi_1
X_1191_ phase_pwm_inst.counter\[18\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0668_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0975_ net88 VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__inv_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1527_ _0490_ net35 _0932_ _0934_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__o221a_1
X_1458_ _0882_ _0883_ _0847_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__and3b_1
X_1389_ _0829_ _0832_ _0830_ _0831_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or4b_1
XFILLER_27_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1174_ phase_pwm_inst.counter\[13\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0651_ sky130_fd_sc_hd__and2_1
X_1312_ _0627_ _0629_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_22_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1243_ _0608_ _0670_ _0671_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__a21boi_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0958_ phase_pwm_inst.counter\[15\] VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__inv_2
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_83 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1930_ clknet_3_5__leaf_clk _0039_ _0113_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 PWM_CNTB[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 PWM_CNTB[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput11 PWM_CNTA[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
Xinput66 TIMER_TOP[10] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
Xinput55 PWM_CNTB[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput22 PWM_CNTA[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput88 TIMER_TOP[30] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
X_1861_ net99 VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__inv_2
Xinput77 TIMER_TOP[20] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
X_1792_ net99 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__inv_2
Xinput99 reset VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_16
X_1226_ _0695_ _0696_ _0616_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__a21oi_1
X_1157_ phase_pwm_inst.counter\[5\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0634_
+ sky130_fd_sc_hd__nor2_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1088_ _0562_ _0563_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1011_ fast_pwm_inst.pwm_counter\[12\] VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__inv_2
X_1913_ clknet_3_1__leaf_clk _0198_ _0096_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[26\]
+ sky130_fd_sc_hd__dfrtp_4
X_1775_ normal_mode_inst.timer_cnt\[25\] _0777_ normal_mode_inst.timer_cnt\[26\] VGND
+ VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a21oi_1
X_1844_ net99 VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_12_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1209_ _0685_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__inv_2
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1560_ fast_pwm_inst.pwm_counter\[14\] _0533_ _0534_ fast_pwm_inst.pwm_counter\[13\]
+ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__o22a_1
X_1491_ fast_pwm_inst.pwm_counter\[30\] _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__or2_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1827_ net99 VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__inv_2
X_1689_ _0353_ _0356_ _0352_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__or3b_1
X_1758_ _0771_ _0410_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__and2b_1
XFILLER_38_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_248 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0991_ net87 VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__inv_2
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1474_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__inv_2
X_1543_ _0475_ net52 net51 _0476_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
X_1612_ _0471_ net25 _0268_ _0281_ _0278_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__o221a_1
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 PWM_CNTA[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
X_1190_ phase_pwm_inst.counter\[19\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0667_ sky130_fd_sc_hd__xor2_1
X_0974_ net89 VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__inv_2
X_1457_ fast_pwm_inst.pwm_counter\[18\] _0880_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__or2_1
X_1526_ fast_pwm_inst.pwm_counter\[10\] _0518_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nand2_1
XFILLER_42_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1388_ net68 _0489_ _0824_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__a21o_1
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1311_ _0759_ phase_pwm_inst.counter\[3\] _0616_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1173_ _0641_ _0642_ _0649_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__and3_1
X_1242_ _0608_ _0670_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nand2_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0957_ phase_pwm_inst.counter\[16\] VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__inv_2
X_1509_ _0915_ _0917_ _0910_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__o21ba_1
XFILLER_46_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1860_ net99 VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__inv_2
Xinput34 PWM_CNTB[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput78 TIMER_TOP[21] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_1
Xinput89 TIMER_TOP[31] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
Xinput23 PWM_CNTA[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput12 PWM_CNTA[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
Xinput67 TIMER_TOP[11] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput45 PWM_CNTB[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
X_1791_ net99 VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__inv_2
Xinput56 PWM_CNTB[30] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1225_ phase_pwm_inst.counter\[30\] _0700_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__xnor2_1
X_1087_ _0444_ net94 net93 _0445_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__o22a_1
X_1156_ _0446_ _0470_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nor2_1
XFILLER_32_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1010_ fast_pwm_inst.pwm_counter\[13\] VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__inv_2
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ net99 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__inv_2
X_1912_ clknet_3_6__leaf_clk _0197_ _0095_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[25\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1774_ normal_mode_inst.timer_cnt\[25\] _0777_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__xor2_1
X_1208_ phase_pwm_inst.counter\[25\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0685_ sky130_fd_sc_hd__nand2_1
XFILLER_27_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1139_ phase_pwm_inst.direction _0600_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__o21ba_4
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _0904_ _0847_ _0903_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__and3b_1
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1826_ net99 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1688_ _0434_ net10 net9 _0435_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a221o_1
X_1757_ normal_mode_inst.timer_cnt\[13\] normal_mode_inst.timer_cnt\[14\] _0769_ normal_mode_inst.timer_cnt\[15\]
+ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a31o_1
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ _0274_ _0279_ _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a21oi_1
X_0990_ net90 VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__inv_2
XFILLER_8_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1473_ fast_pwm_inst.pwm_counter\[24\] fast_pwm_inst.pwm_counter\[23\] fast_pwm_inst.pwm_counter\[22\]
+ _0888_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__and4_1
X_1542_ _0474_ net53 _0502_ fast_pwm_inst.pwm_counter\[27\] VGND VGND VPWR VPWR _0213_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1809_ net99 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0973_ normal_mode_inst.timer_cnt\[0\] VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
X_1456_ fast_pwm_inst.pwm_counter\[18\] fast_pwm_inst.pwm_counter\[17\] fast_pwm_inst.pwm_counter\[16\]
+ _0876_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__and4_1
X_1525_ _0490_ net35 net64 _0492_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__a221o_1
X_1387_ net69 _0488_ _0489_ net68 VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__o22a_1
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1310_ _0630_ _0758_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__xnor2_1
X_1241_ _0710_ phase_pwm_inst.counter\[24\] _0616_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
XFILLER_2_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1172_ _0645_ _0646_ _0648_ _0644_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__and4b_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0956_ phase_pwm_inst.counter\[17\] VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__inv_2
Xoutput100 net100 VGND VGND VPWR VPWR PWM_OUTA sky130_fd_sc_hd__buf_1
X_1508_ _0911_ _0913_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__a21o_1
X_1439_ fast_pwm_inst.pwm_counter\[12\] _0868_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__or2_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 PWM_CNTA[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlymetal6s2s_1
X_1790_ net99 VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
Xinput57 PWM_CNTB[31] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
Xinput46 PWM_CNTB[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput79 TIMER_TOP[22] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput24 PWM_CNTA[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
Xinput35 PWM_CNTB[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
Xinput68 TIMER_TOP[12] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
X_1224_ _0423_ _0695_ _0699_ _0616_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__a211o_1
XFILLER_37_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1086_ net92 _0446_ phase_pwm_inst.counter\[6\] _0467_ VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__o2bb2a_1
X_1155_ _0619_ _0621_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__and3_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1988_ clknet_3_1__leaf_clk _0035_ _0171_ VGND VGND VPWR VPWR phase_pwm_inst.direction
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_7_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1842_ net99 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__inv_2
X_1773_ _0777_ _0416_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__and2b_1
XFILLER_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1911_ clknet_3_3__leaf_clk _0196_ _0094_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[24\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_4_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1207_ phase_pwm_inst.counter\[27\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0684_ sky130_fd_sc_hd__xnor2_1
X_1069_ _0431_ net78 VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1138_ _0606_ _0610_ _0614_ phase_pwm_inst.direction VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__o31a_1
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1756_ normal_mode_inst.timer_cnt\[14\] _0770_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__xnor2_1
X_1825_ net99 VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__inv_2
X_1687_ phase_pwm_inst.counter\[19\] _0528_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1610_ _0269_ _0273_ _0270_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a21bo_1
XFILLER_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1472_ _0891_ _0892_ _0847_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__and3b_1
X_1541_ _0912_ _0208_ _0209_ _0211_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__or4_1
XFILLER_39_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1739_ normal_mode_inst.timer_cnt\[4\] _0763_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__or2_1
X_1808_ net99 VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_2
XFILLER_41_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ phase_pwm_inst.counter\[0\] VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__inv_2
X_1524_ fast_pwm_inst.pwm_counter\[10\] _0518_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_1
X_1455_ _0880_ _0881_ _0847_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__and3b_1
X_1386_ _0465_ fast_pwm_inst.pwm_counter\[11\] _0823_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__nor3_1
XFILLER_50_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1171_ phase_pwm_inst.counter\[11\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0648_ sky130_fd_sc_hd__xor2_1
X_1240_ _0680_ _0691_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0955_ phase_pwm_inst.counter\[18\] VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__inv_2
X_1507_ fast_pwm_inst.pwm_counter\[21\] _0507_ _0508_ fast_pwm_inst.pwm_counter\[20\]
+ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a22o_1
Xoutput101 net101 VGND VGND VPWR VPWR PWM_OUTB sky130_fd_sc_hd__buf_1
X_1369_ net92 _0496_ _0805_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__o22a_1
X_1438_ fast_pwm_inst.pwm_counter\[12\] fast_pwm_inst.pwm_counter\[11\] fast_pwm_inst.pwm_counter\[10\]
+ _0864_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__and4_1
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 PWM_CNTA[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput36 PWM_CNTB[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_1
Xinput14 PWM_CNTA[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput58 PWM_CNTB[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
Xinput47 PWM_CNTB[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput69 TIMER_TOP[13] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1223_ phase_pwm_inst.counter\[29\] _0696_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1154_ _0627_ _0629_ _0622_ _0623_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__a211o_1
X_1085_ _0558_ _0560_ _0561_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a21bo_1
XFILLER_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1987_ clknet_3_6__leaf_clk _0036_ _0170_ VGND VGND VPWR VPWR phase_pwm_inst.pwm_outa
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1910_ clknet_3_2__leaf_clk _0195_ _0093_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[23\]
+ sky130_fd_sc_hd__dfrtp_4
X_1841_ net99 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__inv_2
X_1772_ normal_mode_inst.timer_cnt\[23\] normal_mode_inst.timer_cnt\[22\] _0775_ normal_mode_inst.timer_cnt\[24\]
+ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a31o_1
XFILLER_6_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1137_ _0611_ _0613_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__or2_1
X_1206_ _0681_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__nand2_1
XFILLER_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ _0434_ net74 VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1686_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__inv_2
X_1755_ _0770_ _0409_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_1
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1824_ net99 VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__inv_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _0910_ _0913_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__nand3b_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1471_ _0479_ _0890_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nand2_1
X_1807_ net99 VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_1669_ _0323_ _0337_ _0326_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o21ba_1
X_1738_ _0763_ _0402_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__nor2_1
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0971_ phase_pwm_inst.counter\[1\] VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__inv_2
X_1454_ _0485_ _0878_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__nand2_1
X_1523_ _0492_ net64 net63 _0493_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__o221a_1
X_1385_ _0826_ _0828_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__or2_1
XFILLER_50_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1170_ _0645_ _0646_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__nand2b_1
XFILLER_32_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0954_ phase_pwm_inst.counter\[19\] VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__inv_2
X_1506_ _0914_ _0912_ _0913_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__and3b_1
Xoutput102 net102 VGND VGND VPWR VPWR timer_interrupt sky130_fd_sc_hd__buf_1
X_1437_ _0868_ _0869_ _0847_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__and3b_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1368_ _0809_ _0810_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__a21boi_1
X_1299_ _0638_ _0751_ _0637_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o21ba_1
XFILLER_23_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput26 PWM_CNTA[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput48 PWM_CNTB[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xinput59 PWM_CNTB[4] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 PWM_CNTA[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
Xinput37 PWM_CNTB[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlymetal6s2s_1
X_1222_ phase_pwm_inst.counter\[31\] _0698_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__xnor2_1
X_1084_ _0446_ net92 net91 _0447_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__o22a_1
X_1153_ _0627_ _0629_ _0623_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__a21oi_1
XFILLER_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1986_ clknet_3_6__leaf_clk _0037_ _0169_ VGND VGND VPWR VPWR phase_pwm_inst.pwm_outb
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1840_ net99 VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__inv_2
XFILLER_42_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_1771_ normal_mode_inst.timer_cnt\[23\] _0776_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1067_ _0433_ net75 _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__a21oi_1
X_1136_ phase_pwm_inst.counter\[15\] phase_pwm_inst.counter\[14\] phase_pwm_inst.counter\[13\]
+ phase_pwm_inst.counter\[12\] VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__or4_1
X_1205_ phase_pwm_inst.counter\[26\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0682_ sky130_fd_sc_hd__nand2_1
XFILLER_25_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1969_ clknet_3_0__leaf_clk _0006_ _0152_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1823_ net99 VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__inv_2
X_1685_ phase_pwm_inst.counter\[19\] _0528_ _0529_ phase_pwm_inst.counter\[18\] VGND
+ VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a22o_1
X_1754_ normal_mode_inst.timer_cnt\[13\] _0769_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__or2_1
X_1119_ _0586_ _0591_ _0592_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_0_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1470_ _0479_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_30_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1806_ net99 VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__inv_2
X_1599_ fast_pwm_inst.pwm_counter\[28\] _0521_ _0522_ fast_pwm_inst.pwm_counter\[27\]
+ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a22o_1
X_1668_ _0424_ net53 _0331_ _0335_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o221a_1
X_1737_ normal_mode_inst.timer_cnt\[3\] _0762_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_51_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0970_ phase_pwm_inst.counter\[2\] VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__inv_2
X_1453_ _0485_ _0878_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_1
X_1522_ _0928_ _0929_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a21o_1
XFILLER_4_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1384_ net70 _0487_ _0488_ net69 _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a221o_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0953_ phase_pwm_inst.counter\[20\] VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__inv_2
X_1505_ _0484_ net42 net41 _0485_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__a22o_1
X_1367_ net91 _0497_ _0498_ net90 VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__o22a_1
X_1436_ _0490_ _0866_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__nand2_1
X_1298_ _0633_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nor2_1
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput49 PWM_CNTB[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput16 PWM_CNTA[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 PWM_CNTA[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 PWM_CNTB[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
X_1221_ _0602_ _0696_ _0697_ _0695_ _0616_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a221o_1
X_1083_ phase_pwm_inst.counter\[3\] _0468_ _0557_ _0559_ VGND VGND VPWR VPWR _0560_
+ sky130_fd_sc_hd__a22o_1
X_1152_ _0623_ _0628_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__nor2_1
X_1985_ clknet_3_6__leaf_clk _0024_ _0168_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1419_ _0856_ _0857_ _0847_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__and3b_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1770_ _0776_ _0415_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__and2_1
XFILLER_42_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1204_ phase_pwm_inst.counter\[26\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0681_ sky130_fd_sc_hd__or2_1
X_1066_ _0432_ net77 VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__and2_1
X_1135_ phase_pwm_inst.direction _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__and2_1
X_1899_ clknet_3_0__leaf_clk _0184_ _0082_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_1968_ clknet_3_0__leaf_clk _0005_ _0151_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1753_ _0769_ _0408_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__and2b_1
X_1822_ net99 VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__inv_2
X_1684_ phase_pwm_inst.counter\[17\] _0530_ _0531_ phase_pwm_inst.counter\[16\] VGND
+ VGND VPWR VPWR _0352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1049_ net13 VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__inv_2
X_1118_ _0590_ _0592_ _0594_ _0584_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__and4b_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ _0762_ _0401_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__nor2_1
X_1805_ net99 VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__inv_2
X_1598_ _0471_ net25 net24 _0472_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a22o_1
X_1667_ _0328_ _0329_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
XFILLER_45_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1452_ _0847_ _0878_ _0879_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__and3_1
XFILLER_4_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1521_ _0493_ net63 net62 _0494_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a22o_1
X_1383_ _0463_ fast_pwm_inst.pwm_counter\[15\] VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__nor2_1
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1719_ _0439_ net4 _0385_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__a211o_1
XFILLER_41_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_31 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0952_ phase_pwm_inst.counter\[21\] VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__inv_2
X_1504_ fast_pwm_inst.pwm_counter\[20\] _0508_ _0509_ fast_pwm_inst.pwm_counter\[19\]
+ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__o22a_1
X_1366_ _0468_ fast_pwm_inst.pwm_counter\[3\] fast_pwm_inst.pwm_counter\[2\] _0469_
+ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__o22a_1
X_1435_ _0490_ _0866_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nor2_1
X_1297_ _0634_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__nor2_1
XFILLER_2_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput39 PWM_CNTB[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xinput28 PWM_CNTA[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
Xinput17 PWM_CNTA[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1220_ phase_pwm_inst.counter\[30\] phase_pwm_inst.counter\[29\] VGND VGND VPWR VPWR
+ _0697_ sky130_fd_sc_hd__nand2_1
X_1151_ phase_pwm_inst.counter\[2\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0628_
+ sky130_fd_sc_hd__nor2_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1082_ phase_pwm_inst.counter\[3\] _0468_ _0469_ phase_pwm_inst.counter\[2\] VGND
+ VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o22a_1
X_1984_ clknet_3_7__leaf_clk _0023_ _0167_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[30\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1349_ _0459_ fast_pwm_inst.pwm_counter\[23\] fast_pwm_inst.pwm_counter\[22\] _0460_
+ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__a22o_1
X_1418_ _0496_ _0854_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nand2_1
XFILLER_22_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1134_ phase_pwm_inst.counter\[11\] phase_pwm_inst.counter\[10\] phase_pwm_inst.counter\[9\]
+ phase_pwm_inst.counter\[8\] VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__or4_1
X_1203_ phase_pwm_inst.direction _0610_ _0670_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__o2bb2a_1
X_1065_ phase_pwm_inst.counter\[16\] _0462_ _0540_ _0541_ VGND VGND VPWR VPWR _0542_
+ sky130_fd_sc_hd__a31o_1
X_1898_ clknet_3_0__leaf_clk _0183_ _0081_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_1967_ clknet_3_0__leaf_clk _0004_ _0150_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1683_ _0431_ net14 net13 _0432_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a22o_1
XFILLER_30_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1752_ normal_mode_inst.timer_cnt\[11\] normal_mode_inst.timer_cnt\[10\] _0767_ normal_mode_inst.timer_cnt\[12\]
+ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__a31o_1
X_1821_ net99 VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__inv_2
X_1117_ _0424_ net85 net84 _0425_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__o221a_1
X_1048_ net14 VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1666_ phase_pwm_inst.counter\[25\] _0503_ _0324_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o21ai_1
X_1804_ net99 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_1735_ normal_mode_inst.timer_cnt\[0\] normal_mode_inst.timer_cnt\[1\] normal_mode_inst.timer_cnt\[2\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__a21oi_1
X_1597_ _0251_ _0260_ _0261_ _0266_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__o211a_1
XFILLER_38_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1520_ _0494_ net62 net61 _0495_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__o22a_1
X_1451_ fast_pwm_inst.pwm_counter\[16\] _0876_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__or2_1
X_1382_ net70 _0487_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__o21ai_1
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1649_ _0310_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or2_1
X_1718_ phase_pwm_inst.counter\[13\] _0534_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nor2_1
XFILLER_41_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0951_ phase_pwm_inst.counter\[22\] VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__inv_2
XFILLER_32_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1503_ fast_pwm_inst.pwm_counter\[17\] _0511_ _0512_ fast_pwm_inst.pwm_counter\[16\]
+ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a221o_1
X_1365_ _0469_ fast_pwm_inst.pwm_counter\[2\] _0806_ _0807_ _0808_ VGND VGND VPWR
+ VPWR _0809_ sky130_fd_sc_hd__a221o_1
X_1434_ _0847_ _0866_ _0867_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and3_1
X_1296_ _0617_ _0632_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__nor2_1
XFILLER_11_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 PWM_CNTA[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
Xinput29 PWM_CNTA[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
X_1150_ phase_pwm_inst.counter\[0\] _0625_ _0624_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21bo_1
X_1081_ _0447_ net91 VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__nand2_1
X_1983_ clknet_3_6__leaf_clk _0021_ _0166_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1417_ _0496_ _0854_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__nor2_1
X_1348_ _0459_ fast_pwm_inst.pwm_counter\[23\] VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__nor2_1
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1279_ _0653_ _0732_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_38_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1064_ _0434_ net74 net73 _0435_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__o22ai_1
X_1133_ _0607_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__or2_1
X_1202_ _0673_ _0676_ _0677_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__or3_1
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1966_ clknet_3_1__leaf_clk _0003_ _0149_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_47_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1897_ clknet_3_0__leaf_clk _0182_ _0080_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_34_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1820_ net99 VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__inv_2
X_1682_ _0429_ net16 _0349_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__o21a_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ normal_mode_inst.timer_cnt\[11\] _0768_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_48_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1047_ net17 VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__inv_2
X_1116_ _0422_ net88 net86 _0423_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_0_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1949_ clknet_3_7__leaf_clk _0059_ _0132_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_23_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_8_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1803_ net99 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1596_ _0252_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__or2_1
X_1665_ _0322_ _0327_ _0331_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or4_1
XFILLER_7_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1734_ normal_mode_inst.timer_cnt\[0\] normal_mode_inst.timer_cnt\[1\] VGND VGND
+ VPWR VPWR _0049_ sky130_fd_sc_hd__xor2_1
XFILLER_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1450_ fast_pwm_inst.pwm_counter\[16\] _0876_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__nand2_1
X_1381_ _0463_ fast_pwm_inst.pwm_counter\[15\] VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__nand2_1
XFILLER_50_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1648_ phase_pwm_inst.counter\[18\] _0510_ _0511_ phase_pwm_inst.counter\[17\] _0311_
+ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o221a_1
X_1717_ phase_pwm_inst.counter\[13\] _0534_ _0535_ phase_pwm_inst.counter\[12\] VGND
+ VGND VPWR VPWR _0385_ sky130_fd_sc_hd__a22o_1
X_1579_ _0489_ net4 net3 _0490_ _0228_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__a221o_1
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0950_ phase_pwm_inst.counter\[23\] VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__inv_2
X_1502_ fast_pwm_inst.pwm_counter\[19\] _0509_ _0510_ fast_pwm_inst.pwm_counter\[18\]
+ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a22o_1
X_1433_ fast_pwm_inst.pwm_counter\[10\] _0864_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__or2_1
X_1364_ net76 fast_pwm_inst.pwm_counter\[1\] VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__and2b_1
X_1295_ _0643_ _0748_ phase_pwm_inst.counter\[8\] _0616_ VGND VGND VPWR VPWR _0180_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput19 PWM_CNTA[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ phase_pwm_inst.counter\[2\] _0469_ _0554_ _0555_ _0556_ VGND VGND VPWR VPWR
+ _0557_ sky130_fd_sc_hd__a221o_1
X_1982_ clknet_3_6__leaf_clk _0020_ _0165_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_21_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1347_ _0452_ fast_pwm_inst.pwm_counter\[31\] VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__nor2_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1416_ _0847_ _0854_ _0855_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__and3_1
XFILLER_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1278_ _0737_ phase_pwm_inst.counter\[14\] _0616_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_51_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1201_ _0677_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__inv_2
X_1063_ _0435_ net73 VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_1
X_1132_ phase_pwm_inst.counter\[23\] phase_pwm_inst.counter\[22\] phase_pwm_inst.counter\[21\]
+ phase_pwm_inst.counter\[20\] VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or4_1
XFILLER_33_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1965_ clknet_3_1__leaf_clk _0002_ _0148_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_1896_ clknet_3_0__leaf_clk _0181_ _0079_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1750_ _0768_ _0407_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and2_1
X_1681_ _0429_ net16 net15 _0430_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1046_ net18 VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__inv_2
X_1115_ _0427_ net82 net81 _0428_ _0591_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_0_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1879_ net99 VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
X_1948_ clknet_3_7__leaf_clk _0058_ _0131_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1733_ _0421_ net25 _0339_ _0400_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__o22a_1
X_1802_ net99 VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__inv_2
X_1595_ _0481_ net14 _0254_ _0264_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__o22a_1
X_1664_ _0427_ net50 net49 _0428_ _0332_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a221o_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1029_ net46 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__inv_2
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1380_ net67 _0490_ _0820_ _0822_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__o221a_1
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1716_ _0438_ net6 _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a211o_1
X_1647_ _0308_ _0312_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2b_1
XFILLER_6_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1578_ _0490_ net3 net2 _0491_ _0247_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o221a_1
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1501_ _0480_ net47 net46 _0481_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a22o_1
X_1363_ fast_pwm_inst.pwm_counter\[0\] net65 VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__nand2b_1
X_1432_ fast_pwm_inst.pwm_counter\[10\] _0864_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__nand2_1
XFILLER_48_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1294_ _0641_ _0642_ _0616_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__o21bai_1
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1981_ clknet_3_6__leaf_clk _0019_ _0164_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_15_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1346_ _0781_ _0788_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a21oi_1
XFILLER_28_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1415_ fast_pwm_inst.pwm_counter\[4\] _0852_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1277_ _0654_ _0734_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ phase_pwm_inst.counter\[22\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0677_ sky130_fd_sc_hd__xnor2_2
X_1062_ phase_pwm_inst.counter\[22\] _0460_ _0461_ phase_pwm_inst.counter\[21\] VGND
+ VGND VPWR VPWR _0539_ sky130_fd_sc_hd__o22a_1
X_1131_ phase_pwm_inst.direction _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nand2_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1895_ clknet_3_0__leaf_clk _0180_ _0078_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_1964_ clknet_3_1__leaf_clk _0001_ _0147_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_1329_ normal_mode_inst.timer_cnt\[19\] _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1680_ _0341_ _0347_ _0340_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_48_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1114_ phase_pwm_inst.counter\[26\] _0457_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1045_ net19 VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__inv_2
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1947_ clknet_3_6__leaf_clk _0057_ _0130_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[27\]
+ sky130_fd_sc_hd__dfrtp_1
X_1878_ net99 VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__inv_2
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1663_ _0424_ net53 VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__nor2_1
X_1732_ _0395_ _0396_ _0399_ _0348_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__o31a_1
X_1801_ net99 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__inv_2
X_1594_ _0482_ net13 net11 _0483_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1028_ net47 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__inv_2
XFILLER_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1646_ _0307_ _0309_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__nor3_1
X_1715_ phase_pwm_inst.counter\[15\] _0532_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nor2_1
X_1577_ _0244_ _0245_ _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a21o_1
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1500_ fast_pwm_inst.pwm_counter\[23\] _0505_ _0506_ fast_pwm_inst.pwm_counter\[22\]
+ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a22o_1
X_1293_ _0747_ phase_pwm_inst.counter\[9\] _0616_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
X_1362_ fast_pwm_inst.pwm_counter\[1\] net76 VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__nand2b_1
X_1431_ _0864_ _0865_ _0847_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__and3b_1
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1629_ _0295_ _0296_ _0297_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__a21o_1
XFILLER_45_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1980_ clknet_3_6__leaf_clk _0018_ _0163_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_9_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1345_ _0452_ fast_pwm_inst.pwm_counter\[31\] fast_pwm_inst.pwm_counter\[30\] _0453_
+ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__a22o_1
X_1414_ fast_pwm_inst.pwm_counter\[4\] _0852_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__nand2_1
X_1276_ _0736_ phase_pwm_inst.counter\[15\] _0616_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_51_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1130_ phase_pwm_inst.counter\[19\] phase_pwm_inst.counter\[18\] phase_pwm_inst.counter\[17\]
+ phase_pwm_inst.counter\[16\] VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or4_1
XFILLER_26_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1061_ phase_pwm_inst.counter\[23\] _0459_ _0460_ phase_pwm_inst.counter\[22\] VGND
+ VGND VPWR VPWR _0538_ sky130_fd_sc_hd__a22o_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1963_ clknet_3_0__leaf_clk _0031_ _0146_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_1894_ clknet_3_1__leaf_clk _0179_ _0077_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_1328_ normal_mode_inst.timer_cnt\[17\] normal_mode_inst.timer_cnt\[16\] normal_mode_inst.timer_cnt\[18\]
+ _0771_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_3_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1259_ _0660_ _0662_ _0663_ _0664_ _0668_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__a311oi_1
XTAP_TAPCELL_ROW_34_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1044_ net20 VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__inv_2
X_1113_ _0587_ _0588_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_0_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1877_ net99 VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__inv_2
X_1946_ clknet_3_7__leaf_clk _0056_ _0129_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1800_ net99 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__inv_2
X_1731_ phase_pwm_inst.counter\[24\] _0525_ _0397_ _0398_ VGND VGND VPWR VPWR _0399_
+ sky130_fd_sc_hd__a211o_1
X_1662_ _0328_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__nand2_1
X_1593_ _0253_ _0262_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__or2_1
X_1027_ net48 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__inv_2
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1929_ clknet_3_5__leaf_clk _0069_ _0112_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1645_ _0310_ _0311_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or3_1
X_1576_ _0491_ net2 net32 _0492_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a22o_1
X_1714_ phase_pwm_inst.counter\[14\] _0533_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__a21o_1
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1430_ fast_pwm_inst.pwm_counter\[9\] _0862_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__or2_1
X_1292_ _0647_ _0741_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__xnor2_1
X_1361_ net91 _0497_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__and2_1
X_1628_ _0441_ net34 net64 _0442_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__a22o_1
X_1559_ fast_pwm_inst.pwm_counter\[15\] _0532_ _0533_ fast_pwm_inst.pwm_counter\[14\]
+ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a22o_1
XFILLER_39_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1413_ _0852_ _0853_ _0847_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__and3b_1
X_1344_ _0454_ fast_pwm_inst.pwm_counter\[29\] fast_pwm_inst.pwm_counter\[28\] _0455_
+ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a221o_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1275_ _0656_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__xnor2_1
XFILLER_51_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1060_ _0429_ net80 VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_25_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ clknet_3_1__leaf_clk _0030_ _0145_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_1893_ clknet_3_4__leaf_clk _0178_ _0076_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1327_ normal_mode_inst.timer_cnt\[16\] _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__nand2_1
X_1258_ _0665_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nand2_1
X_1189_ _0663_ _0665_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1043_ net21 VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__inv_2
X_1112_ phase_pwm_inst.counter\[27\] _0456_ _0457_ phase_pwm_inst.counter\[26\] VGND
+ VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1945_ clknet_3_7__leaf_clk _0055_ _0128_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1876_ net99 VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__inv_2
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1592_ _0255_ _0256_ _0484_ net10 VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__o2bb2a_1
X_1661_ _0426_ net51 _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__a21oi_1
X_1730_ _0423_ net22 net21 _0424_ _0343_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a221o_1
XFILLER_11_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1026_ net49 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_28_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1859_ net99 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_12_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1928_ clknet_3_5__leaf_clk _0068_ _0111_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1713_ _0437_ net7 VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__nor2_1
X_1644_ _0436_ net40 net39 _0437_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__a221o_1
X_1575_ _0492_ net32 net31 _0493_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o22a_1
X_1009_ fast_pwm_inst.pwm_counter\[14\] VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__inv_2
XFILLER_25_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1360_ _0794_ _0803_ _0793_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1291_ _0746_ phase_pwm_inst.counter\[10\] _0616_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_16_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1489_ fast_pwm_inst.pwm_counter\[29\] fast_pwm_inst.pwm_counter\[28\] _0900_ VGND
+ VGND VPWR VPWR _0904_ sky130_fd_sc_hd__and3_1
X_1627_ _0442_ net64 net63 _0443_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__o22a_1
X_1558_ fast_pwm_inst.pwm_counter\[15\] _0532_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__nor2_1
XFILLER_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1343_ _0455_ fast_pwm_inst.pwm_counter\[28\] _0785_ _0786_ VGND VGND VPWR VPWR _0787_
+ sky130_fd_sc_hd__o22a_1
X_1412_ fast_pwm_inst.pwm_counter\[3\] _0851_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__or2_1
XFILLER_36_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1274_ _0652_ _0654_ _0733_ phase_pwm_inst.direction phase_pwm_inst.counter\[14\]
+ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__a32o_1
X_0989_ net93 VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__inv_2
XFILLER_42_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1961_ clknet_3_1__leaf_clk _0029_ _0144_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_18_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1892_ clknet_3_1__leaf_clk _0177_ _0075_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1326_ normal_mode_inst.timer_cnt\[13\] normal_mode_inst.timer_cnt\[15\] normal_mode_inst.timer_cnt\[14\]
+ _0769_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_3_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1188_ phase_pwm_inst.counter\[17\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0665_ sky130_fd_sc_hd__or2_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1257_ _0660_ _0662_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_42_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1042_ net22 VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__inv_2
X_1111_ _0421_ net89 net88 _0422_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1875_ net99 VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__inv_2
X_1944_ clknet_3_7__leaf_clk _0054_ _0127_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1309_ _0620_ _0622_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_22_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1591_ _0479_ net16 net15 _0480_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o22a_1
X_1660_ phase_pwm_inst.counter\[27\] _0502_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nor2_1
XFILLER_7_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1025_ net50 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__inv_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1858_ net99 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__inv_2
X_1927_ clknet_3_5__leaf_clk _0067_ _0110_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1789_ net99 VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__inv_2
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1643_ phase_pwm_inst.counter\[23\] _0505_ _0506_ phase_pwm_inst.counter\[22\] VGND
+ VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a22o_1
XANTENNA_1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1712_ _0374_ _0377_ _0379_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__o21a_1
XFILLER_6_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1574_ _0241_ _0242_ _0243_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a21o_1
X_1008_ fast_pwm_inst.pwm_counter\[16\] VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__inv_2
XFILLER_32_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1290_ _0644_ _0742_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__xnor2_1
XFILLER_31_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1626_ _0292_ _0293_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a21o_1
X_1488_ _0473_ _0902_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nand2_1
X_1557_ _0215_ _0218_ _0223_ _0227_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o211a_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1342_ net84 _0475_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__nor2_1
X_1411_ fast_pwm_inst.pwm_counter\[3\] fast_pwm_inst.pwm_counter\[2\] fast_pwm_inst.pwm_counter\[1\]
+ fast_pwm_inst.pwm_counter\[0\] VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__and4_1
X_1273_ _0652_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__nand2_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0988_ net95 VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1609_ fast_pwm_inst.pwm_counter\[26\] _0523_ _0271_ _0276_ VGND VGND VPWR VPWR _0279_
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1960_ clknet_3_1__leaf_clk _0028_ _0143_ VGND VGND VPWR VPWR fast_pwm_inst.pwm_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_1891_ clknet_3_4__leaf_clk _0176_ _0074_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1325_ normal_mode_inst.timer_cnt\[13\] _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nand2_1
X_1256_ _0721_ phase_pwm_inst.counter\[20\] _0616_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
X_1187_ phase_pwm_inst.counter\[17\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0664_ sky130_fd_sc_hd__nor2_1
X_1110_ _0428_ net81 _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__a211o_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1041_ net58 VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__inv_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1874_ net99 VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__inv_2
X_1943_ clknet_3_7__leaf_clk _0053_ _0126_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1239_ _0709_ phase_pwm_inst.counter\[25\] _0616_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
X_1308_ _0757_ phase_pwm_inst.counter\[4\] _0616_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1590_ fast_pwm_inst.pwm_counter\[18\] _0529_ net9 _0485_ _0259_ VGND VGND VPWR VPWR
+ _0260_ sky130_fd_sc_hd__a221o_1
XFILLER_7_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1024_ net52 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__inv_2
X_1857_ net99 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__inv_2
X_1788_ net99 VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__inv_2
X_1926_ clknet_3_5__leaf_clk _0066_ _0109_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1642_ phase_pwm_inst.counter\[17\] _0511_ _0512_ phase_pwm_inst.counter\[16\] VGND
+ VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a22o_1
X_1711_ _0440_ net3 _0378_ _0441_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o22a_1
X_1573_ _0493_ net31 net30 _0494_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__a22o_1
X_1007_ fast_pwm_inst.pwm_counter\[17\] VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__inv_2
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1909_ clknet_3_3__leaf_clk _0194_ _0092_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1556_ _0471_ net57 _0219_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o22a_1
X_1625_ _0443_ net63 net62 _0444_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a22o_1
X_1487_ _0847_ _0901_ _0902_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__and3_1
XFILLER_36_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ _0851_ _0847_ _0850_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__and3b_1
X_1341_ _0783_ _0784_ _0782_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o21a_1
X_1272_ _0651_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__or2_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0987_ net67 VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1608_ _0267_ _0271_ _0272_ _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__or4b_1
X_1539_ _0914_ _0916_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nor2_1
XFILLER_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1890_ clknet_3_4__leaf_clk _0175_ _0073_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1186_ phase_pwm_inst.counter\[17\] phase_pwm_inst.direction VGND VGND VPWR VPWR
+ _0663_ sky130_fd_sc_hd__nand2_1
X_1324_ normal_mode_inst.timer_cnt\[11\] normal_mode_inst.timer_cnt\[10\] normal_mode_inst.timer_cnt\[12\]
+ _0767_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__and4_1
X_1255_ _0671_ _0711_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1040_ net34 VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__inv_2
X_1942_ clknet_3_7__leaf_clk _0052_ _0125_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1873_ net99 VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1238_ _0688_ _0703_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__xnor2_1
X_1169_ phase_pwm_inst.counter\[9\] phase_pwm_inst.direction VGND VGND VPWR VPWR _0646_
+ sky130_fd_sc_hd__or2_1
X_1307_ _0632_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2b_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_45_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1023_ fast_pwm_inst.pwm_counter\[0\] VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__inv_2
X_1925_ clknet_3_5__leaf_clk _0065_ _0108_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_1856_ net99 VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__inv_2
X_1787_ net99 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1641_ phase_pwm_inst.counter\[19\] _0509_ _0510_ phase_pwm_inst.counter\[18\] VGND
+ VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a22o_1
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1572_ _0494_ net30 net29 _0495_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__o22a_1
X_1710_ net2 _0376_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1006_ fast_pwm_inst.pwm_counter\[18\] VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__inv_2
X_1839_ net99 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__inv_2
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1908_ clknet_3_3__leaf_clk _0193_ _0091_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1555_ _0213_ _0225_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__nor2_1
X_1624_ _0444_ net62 net61 _0445_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__o22a_1
X_1486_ fast_pwm_inst.pwm_counter\[28\] _0900_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__nand2_1
XFILLER_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1340_ net82 _0477_ _0478_ net81 VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__a211oi_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1271_ phase_pwm_inst.counter\[12\] phase_pwm_inst.direction _0731_ VGND VGND VPWR
+ VPWR _0732_ sky130_fd_sc_hd__a21o_1
XFILLER_8_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ net69 VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1469_ fast_pwm_inst.pwm_counter\[22\] _0888_ _0890_ _0847_ VGND VGND VPWR VPWR _0014_
+ sky130_fd_sc_hd__o211a_1
X_1607_ _0476_ net19 _0274_ _0275_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__o2111a_1
X_1538_ _0479_ net48 net40 _0486_ _0909_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_6_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1323_ normal_mode_inst.timer_cnt\[10\] _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__nand2_1
XFILLER_5_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1254_ _0720_ phase_pwm_inst.counter\[21\] _0616_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
X_1185_ _0661_ _0658_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__nand2b_1
XFILLER_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ phase_pwm_inst.counter\[3\] VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_2_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1872_ net99 VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__inv_2
X_1941_ clknet_3_7__leaf_clk _0051_ _0124_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_1306_ _0621_ _0631_ _0619_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_46_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1168_ _0442_ _0470_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__nor2_1
X_1099_ _0553_ _0567_ _0568_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__nor3_1
X_1237_ _0708_ phase_pwm_inst.counter\[26\] _0616_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
XFILLER_20_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1022_ fast_pwm_inst.pwm_counter\[1\] VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__inv_2
X_1855_ net99 VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__inv_2
X_1924_ clknet_3_5__leaf_clk _0064_ _0107_ VGND VGND VPWR VPWR normal_mode_inst.timer_cnt\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1786_ net99 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1640_ _0430_ net47 net46 _0431_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a221o_1
XFILLER_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1571_ _0238_ _0240_ _0239_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__a21o_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ fast_pwm_inst.pwm_counter\[19\] VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__inv_2
XFILLER_34_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1838_ net99 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__inv_2
X_1907_ clknet_3_2__leaf_clk _0192_ _0090_ VGND VGND VPWR VPWR phase_pwm_inst.counter\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_1769_ normal_mode_inst.timer_cnt\[22\] _0775_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__or2_1
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_33_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1485_ fast_pwm_inst.pwm_counter\[28\] _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__or2_1
XFILLER_39_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1554_ _0220_ _0224_ _0214_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a21oi_1
X_1623_ _0445_ net61 _0284_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a22o_1
.ends

